* Component: $AnalogIP/default.group/logic.views/testBuffer  Viewpoint: eldonet
.INCLUDE $AnalogIP/default.group/logic.views/testBuffer/eldonet/testBuffer_eldonet.spi
.INCLUDE $MGC_DESIGN_KIT/models/ELDO/include_all
.PROBE VX




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 
.PARAM Ib=20u 
.STEP PARAM  Ib 20u 60u LIN 10 

.AC dec 10 1 10gig

