*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Mon Nov  4 2013 at 13:54:58

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/folded
*
        M29 VB2T VB2T N$539 VDD p_33_mm l=1u w=14u ad=8.96p as=8.96p pd=29.28u
+  ps=29.28u m=1
        M3 N$431 CMFB VDD VDD p_33_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*8.4e-07)/2):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*6.4e-07+(1-2)/2*({(Wl/1)}*8.4e-07))/1):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+8.4e-07):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+6.4e-07)+(1-2)*({(Wl/1)}+8.4e-07))/1):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  m=1
        C6 VI- VO+ 1P
        M1 N$434 VI+ N$531 VDD p_33_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*8.4e-07)/2):(({(Win/1)}*6.4e-07+((1-1)*{(Win/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*6.4e-07+(1-2)/2*({(Win/1)}*8.4e-07))/1):(({(Win/1)}*6.4e-07+((1-1)*{(Win/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+8.4e-07):((2*({(Win/1)}+6.4e-07)+(1-1)*({(Win/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+6.4e-07)+(1-2)*({(Win/1)}+8.4e-07))/1):((2*({(Win/1)}+6.4e-07)+(1-1)*({(Win/1)}+8.4e-07))/1))}
+  m=1
        M7 N$437 VB4 GROUND GROUND n_33_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*8.4e-07)/2):(({(Wf/1)}*6.4e-07+((1-1)*{(Wf/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*6.4e-07+(1-2)/2*({(Wf/1)}*8.4e-07))/1):(({(Wf/1)}*6.4e-07+((1-1)*{(Wf/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+8.4e-07):((2*({(Wf/1)}+6.4e-07)+(1-1)*({(Wf/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+6.4e-07)+(1-2)*({(Wf/1)}+8.4e-07))/1):((2*({(Wf/1)}+6.4e-07)+(1-1)*({(Wf/1)}+8.4e-07))/1))}
+  m=1
        M4 VO- VB2 N$431 VDD p_33_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*8.4e-07)/2):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*6.4e-07+(1-2)/2*({(Wcl/1)}*8.4e-07))/1):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+8.4e-07):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+6.4e-07)+(1-2)*({(Wcl/1)}+8.4e-07))/1):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  m=1
        M8 N$434 VB4 GROUND GROUND n_33_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*8.4e-07)/2):(({(Wf/1)}*6.4e-07+((1-1)*{(Wf/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*6.4e-07+(1-2)/2*({(Wf/1)}*8.4e-07))/1):(({(Wf/1)}*6.4e-07+((1-1)*{(Wf/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+8.4e-07):((2*({(Wf/1)}+6.4e-07)+(1-1)*({(Wf/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+6.4e-07)+(1-2)*({(Wf/1)}+8.4e-07))/1):((2*({(Wf/1)}+6.4e-07)+(1-1)*({(Wf/1)}+8.4e-07))/1))}
+  m=1
        E3 N$493 GROUND Vo- 0 0.5
        E2 N$494 N$493 Vo+ 0 0.5
        E5 VDD CMFB N$494 VOCM -10
        M25 N$531 VB2T N$532 VDD p_33_mm l=1u w=100u ad=64p as=64p pd=0.201m
+  ps=0.201m m=1
        M32 VB4 VB4 GROUND GROUND n_33_mm l=Lf w={{({Wf/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wf/2}/1)}*8.4e-07)/2):(({({Wf/2}/1)}*6.4e-07+((1-1)*{({Wf/2}/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wf/2}/1)}*6.4e-07+(1-2)/2*({({Wf/2}/1)}*8.4e-07))/1):(({({Wf/2}/1)}*6.4e-07+((1-1)*{({Wf/2}/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wf/2}/1)}+8.4e-07):((2*({({Wf/2}/1)}+6.4e-07)+(1-1)*({({Wf/2}/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wf/2}/1)}+6.4e-07)+(1-2)*({({Wf/2}/1)}+8.4e-07))/1):((2*({({Wf/2}/1)}+6.4e-07)+(1-1)*({({Wf/2}/1)}+8.4e-07))/1))}
+  m=1
        M33 VB3 VB3 VB4 GROUND n_33_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*8.4e-07)/2):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*6.4e-07+(1-2)/2*({(Wcf/1)}*8.4e-07))/1):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+8.4e-07):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+6.4e-07)+(1-2)*({(Wcf/1)}+8.4e-07))/1):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  m=1
        M20 VO- VB3 N$434 GROUND n_33_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*8.4e-07)/2):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*6.4e-07+(1-2)/2*({(Wcf/1)}*8.4e-07))/1):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+8.4e-07):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+6.4e-07)+(1-2)*({(Wcf/1)}+8.4e-07))/1):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  m=1
        C3 VOCM VO- 0.5P
        E4 VO GROUND VO- VO+ 1
        M31 N$571 N$571 VDD VDD p_33_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*8.4e-07)/2):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*6.4e-07+(1-2)/2*({(Wl/1)}*8.4e-07))/1):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+8.4e-07):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+6.4e-07)+(1-2)*({(Wl/1)}+8.4e-07))/1):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  m=1
        C5 VI+ VO- 1P
        M30 VB2 VB2 N$571 VDD p_33_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*8.4e-07)/2):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*6.4e-07+(1-2)/2*({(Wcl/1)}*8.4e-07))/1):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+8.4e-07):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+6.4e-07)+(1-2)*({(Wcl/1)}+8.4e-07))/1):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  m=1
        M6 VO+ VB2 N$433 VDD p_33_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*8.4e-07)/2):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*6.4e-07+(1-2)/2*({(Wcl/1)}*8.4e-07))/1):(({(Wcl/1)}*6.4e-07+((1-1)*{(Wcl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+8.4e-07):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+6.4e-07)+(1-2)*({(Wcl/1)}+8.4e-07))/1):((2*({(Wcl/1)}+6.4e-07)+(1-1)*({(Wcl/1)}+8.4e-07))/1))}
+  m=1
        M2 N$437 VI- N$531 VDD p_33_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*8.4e-07)/2):(({(Win/1)}*6.4e-07+((1-1)*{(Win/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*6.4e-07+(1-2)/2*({(Win/1)}*8.4e-07))/1):(({(Win/1)}*6.4e-07+((1-1)*{(Win/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+8.4e-07):((2*({(Win/1)}+6.4e-07)+(1-1)*({(Win/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+6.4e-07)+(1-2)*({(Win/1)}+8.4e-07))/1):((2*({(Win/1)}+6.4e-07)+(1-1)*({(Win/1)}+8.4e-07))/1))}
+  m=1
        R4 N$579 VI+ 100gig
        R3 N$584 VI- 100gig
        V1 N$575 GROUND PULSE ( 0V 0.1V 10nS 0.01nS 0.01nS 15nS 30nS )
        R1 VI+ VO- 100gig
        R2 VI- VO+ 100gig
        V3 VDD GROUND DC 3.3V
        C7 N$584 VI- 0.25P
        I4 VB2 VB3 DC 70u
        V2 VOCM GROUND DC 1.6
        C2 N$579 VI+ 0.25P
        C4 VO+ VOCM 0.5P
        M9 VO+ VB3 N$437 GROUND n_33_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*8.4e-07)/2):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*6.4e-07+(1-2)/2*({(Wcf/1)}*8.4e-07))/1):(({(Wcf/1)}*6.4e-07+((1-1)*{(Wcf/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+8.4e-07):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+6.4e-07)+(1-2)*({(Wcf/1)}+8.4e-07))/1):((2*({(Wcf/1)}+6.4e-07)+(1-1)*({(Wcf/1)}+8.4e-07))/1))}
+  m=1
        M24 N$532 VB1T VDD VDD p_33_mm l=1u w=100u ad=64p as=64p pd=0.201m
+  ps=0.201m m=1
        M5 N$433 CMFB VDD VDD p_33_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*8.4e-07)/2):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*6.4e-07+(1-2)/2*({(Wl/1)}*8.4e-07))/1):(({(Wl/1)}*6.4e-07+((1-1)*{(Wl/1)}*8.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+8.4e-07):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+6.4e-07)+(1-2)*({(Wl/1)}+8.4e-07))/1):((2*({(Wl/1)}+6.4e-07)+(1-1)*({(Wl/1)}+8.4e-07))/1))}
+  m=1
        V6 N$478 GROUND DC 1.6
        X_S2D2 N$579 N$584 N$478 N$575 GROUND S2D
        M28 N$529 VB1T VDD VDD p_33_mm l=1u w=14u ad=8.96p as=8.96p pd=29.28u
+  ps=29.28u m=1
        M27 VB1T VB2T N$529 VDD p_33_mm l=1u w=14u ad=8.96p as=8.96p pd=29.28u
+  ps=29.28u m=1
        M26 N$539 VB2T VDD VDD p_33_mm l=5u w=14u ad=8.96p as=8.96p pd=29.28u
+  ps=29.28u m=1
        I3 VB1T GROUND DC 20u
        I2 VB2T GROUND DC 20u
*
.end
