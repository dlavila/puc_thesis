*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Thu Jan  9 2014 at 13:27:18

*
* Globals.
*
.global VDD GROUND


*
* Component pathname : $MGC_DESIGN_KIT/symbols/RNHR1000_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/RNHR1000_MM/rnhr1000_mm


*
* Component pathname : $MGC_DESIGN_KIT/symbols/MIMCAPS_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/MIMCAPS_MM/mimcaps_mm

*
* Component pathname : $SC_filter/default.group/logic.views/BUFFER
*
.subckt BUFFER  VO AGND AVDD IB VI+ VI-

        M50 N$427 N$427 N$204 AGND n_18_mm l=0.45u w=5.12u ad=1.382p as=1.608p
+  pd=5.66u ps=6.772u m=10
        M45 VB3 IB AVDD AVDD p_18_mm l=0.45u w=5u ad=1.35p as=1.9p pd=5.54u
+  ps=8.26u m=4
        M21 VB3 VB3 N$148 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M24 N$148 VB3 AGND AGND n_18_mm l=2.25u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M49 ND4 N$626 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M47 ND3 N$698 ND3 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M57 ND1 N$681 ND1 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M46 ND4 N$618 ND4 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M44 ND3 N$684 ND3 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        MIN1 ND1 VI- N$204 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.52p
+  pd=2.14u ps=2.65u m=8
        M2 N$165 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p
+  pd=2.14u ps=3.16u m=4
        M8 ND8 VNCAS ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M42 N$427 N$427 N$209 AVDD p_18_mm l=0.45u w=8u ad=2.16p as=2.512p
+  pd=8.54u ps=10.228u m=10
        M33 VPCAS VPCAS N$131 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        XC2 N$356 VO mimcaps_mm w=11u l=11u m=4
        M19 N$427 N$427 N$209 AVDD p_18_mm l=0.45u w=8u ad=2.16p as=2.512p
+  pd=8.54u ps=10.228u m=10
        M15 ND3 ND6 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        M29 N$250 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M7 ND7 VB3 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p pd=2.14u
+  ps=3.16u m=4
        XC1 N$593 VO mimcaps_mm w=11u l=11u m=4
        XR2 ND7 N$593 AGND rnhr1000_mm lr=10u wr=4u m=1
        M12 ND9 VB2 ND2 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M64 ND2 N$671 ND2 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M63 ND1 N$668 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M62 ND4 N$701 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M61 ND3 N$665 ND3 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M56 ND9 N$650 ND9 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M55 ND8 N$695 ND8 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M54 ND7 N$642 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M25 N$247 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M14 ND7 VPCAS ND9 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M27 N$249 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M26 VPCAS VB3 N$249 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M31 N$253 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M76 ND4 N$741 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M75 ND4 N$737 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M68 ND9 N$692 ND9 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M67 ND8 N$676 ND8 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M66 ND7 N$702 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M65 ND6 N$672 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M28 VB2 VB3 N$250 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M3 N$206 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M17 ND2 VI+ N$204 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.52p
+  pd=2.14u ps=2.65u m=8
        M6 ND2 ND8 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p pd=3.04u
+  ps=4.51u m=4
        XR1 ND9 N$356 AGND rnhr1000_mm lr=10u wr=4u m=1
        MOUTN VO ND7 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.467p
+  pd=2.14u ps=2.344u m=20
        M53 ND6 N$696 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M52 ND2 N$689 ND2 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M1 N$209 VB2 N$206 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M11 ND9 VNCAS ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M40 VB1 VB2 N$277 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M18 ND3 VI- N$209 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.744p
+  pd=3.04u ps=3.408u m=16
        M39 VNCAS VB2 N$274 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M74 VB3 N$734 VB3 AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M73 VB3 N$733 VB3 AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M20 ND2 N$683 ND2 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M_D1 ND1 N$610 ND1 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M35 N$255 N$255 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        M43 VB4 IB AVDD AVDD p_18_mm l=0.45u w=5u ad=1.35p as=1.9p pd=5.54u
+  ps=8.26u m=4
        M48 IB IB AVDD AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M4 N$204 VB3 N$165 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p
+  pd=2.14u ps=3.16u m=4
        M10 ND8 VB2 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M34 N$131 N$131 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p
+  pd=3.04u ps=4.51u m=4
        M51 ND1 N$688 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M41 ND4 VI+ N$209 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.744p
+  pd=3.04u ps=3.408u m=16
        M30 VB1 VB3 N$253 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        MOUTP VO ND9 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.702p
+  pd=3.04u ps=3.187u m=40
        M23 VB4 VB3 N$247 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M22 VB2 VB2 N$279 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M38 N$277 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M72 ND4 N$715 ND4 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M71 ND3 N$711 ND3 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M9 ND6 VB3 ND3 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p pd=2.14u
+  ps=3.16u m=4
        M16 ND4 ND6 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        M36 N$279 VB2 AVDD AVDD p_18_mm l=2.25u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M13 ND6 VPCAS ND8 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M60 ND4 N$687 ND4 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M59 ND3 N$660 ND3 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M58 ND2 N$659 ND2 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M32 VNCAS VNCAS N$255 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M70 ND4 N$708 ND4 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M69 ND3 N$705 ND3 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M5 ND1 ND8 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p pd=3.04u
+  ps=4.51u m=4
        M37 N$274 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
.ends BUFFER

*
* MAIN CELL: Component pathname : $SC_filter/default.group/logic.views/testBuffer
*
        V3 N$31 N$29 PULSE ( 0V 1V 10nS 1nS 1nS 200nS 400nS )
        V2 N$29 GROUND DC 0.2V
        C1 VO GROUND 4P
        V1 VDD GROUND DC 1.8V
        I1 N$2 GROUND DC 3.75uA
        X_BUFFER1 VO GROUND VDD N$2 N$31 VO BUFFER
*
.end
