*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Mon Dec 16 2013 at 14:58:08

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $SC_filter/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $LS_BUFFER/default.group/logic.views/NEW_BUFFER
*
        E1 VO GROUND VO+ VO- 1
        C2 VO- GROUND 0.5P
        M6 N$488 N$488 N$489 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M15 N$492 N$489 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M18 N$500 N$501 N$502 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M17 N$502 N$499 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M14 N$501 N$501 N$499 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        I2 N$501 GROUND DC Ib
        M13 N$499 N$499 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M12 N$500 N$500 GROUND GROUND n_18_mm l=Ln w={{({Wn/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/5}/1)}*5.4e-07)/2):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/5}/1)}*4.9e-07+(1-2)/2*({({Wn/5}/1)}*5.4e-07))/1):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/5}/1)}+5.4e-07):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/5}/1)}+4.9e-07)+(1-2)*({({Wn/5}/1)}+5.4e-07))/1):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  m=1
        M16 N$491 N$488 N$492 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M11 N$494 N$500 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M10 VO+ N$499 VDD VDD p_18_mm l=Lp w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        C1 VO+ GROUND 0.5P
        M9 VO+ N$494 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M8 N$494 VI+ VO+ VO+ p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        C6 VO+ N$494 0.1P
        C5 VO- N$453 0.1P
        V3 VDD GROUND DC 1.8V
        V1 N$72 GROUND PULSE ( -0.6V 0.6V 10nS 0.01nS 0.01nS 20nS 40nS )
        I1 N$488 GROUND DC Ib
        M7 N$489 N$489 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M5 N$491 N$491 GROUND GROUND n_18_mm l=Ln w={{({Wn/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/5}/1)}*5.4e-07)/2):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/5}/1)}*4.9e-07+(1-2)/2*({({Wn/5}/1)}*5.4e-07))/1):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/5}/1)}+5.4e-07):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/5}/1)}+4.9e-07)+(1-2)*({({Wn/5}/1)}+5.4e-07))/1):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  m=1
        M2 N$453 N$491 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M1 VO- N$489 VDD VDD p_18_mm l=Lp w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M3 N$453 VI- VO- VO- p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M4 VO- N$453 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        X_S2D1 VI+ VI- N$74 N$72 GROUND S2D
        V2 N$74 GROUND DC 1V
*
.end
