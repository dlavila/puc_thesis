* Component: $AnalogIP/default.group/logic.views/testRFC  Viewpoint: eldonet
.INCLUDE $AnalogIP/default.group/logic.views/testRFC/eldonet/testRFC_eldonet.spi
.INCLUDE $MGC_DESIGN_KIT/models/ELDO/include_all
.PROBE VX
.PROBE I
.PROBE ISUB




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 
.PARAM Ln=0.18u 
.PARAM Vicm=0.7 

.OPTION PROBOP2
.OPTION PROBOPX
.OP
.TRAN  0 200n 0 10p
