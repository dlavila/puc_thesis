*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Wed Nov  6 2013 at 16:53:20

*
* Globals.
*
.global GROUND

*
* Component pathname : $SC_filter/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $SC_filter/default.group/logic.views/RFC3
*
        M14 N$105 VI+ N$23 N$23 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M24 N$195 N$195 GROUND GROUND n_18_mm l=0.5u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        C3 VOCM VO- 1P
        M9 N$17 CMFB VDD VDD p_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        V6 N$28 GROUND DC Vicm
        C2 N$26 VI+ 0.25P
        E4 VO GROUND VO- VO+ 1
        M11 N$98 VB3 N$47 GROUND n_18_mm l=Laux w={{(Waux/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Waux/1)}*5.4e-07)/2):(({(Waux/1)}*4.9e-07+((1-1)*{(Waux/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Waux/1)}*4.9e-07+(1-2)/2*({(Waux/1)}*5.4e-07))/1):(({(Waux/1)}*4.9e-07+((1-1)*{(Waux/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Waux/1)}+5.4e-07):((2*({(Waux/1)}+4.9e-07)+(1-1)*({(Waux/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Waux/1)}+4.9e-07)+(1-2)*({(Waux/1)}+5.4e-07))/1):((2*({(Waux/1)}+4.9e-07)+(1-1)*({(Waux/1)}+5.4e-07))/1))}
+  m=1
        X_S2D2 N$26 N$124 N$28 N$29 GROUND S2D
        M10 N$101 CMFB VDD VDD p_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        C4 VO+ VOCM 1P
        M2 VB1T VB1T VDD VDD p_18_mm l=0.5u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        E6 N$41 GROUND Vo- 0 0.5
        M8 VO+ VB2 N$101 VDD p_18_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*5.4e-07)/2):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*4.9e-07+(1-2)/2*({(Wcl/1)}*5.4e-07))/1):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+5.4e-07):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+4.9e-07)+(1-2)*({(Wcl/1)}+5.4e-07))/1):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  m=1
        C5 VI+ VO- 1P
        M5 VO- VB3 N$5 GROUND n_18_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*5.4e-07)/2):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*4.9e-07+(1-2)/2*({(Wcf/1)}*5.4e-07))/1):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+5.4e-07):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+4.9e-07)+(1-2)*({(Wcf/1)}+5.4e-07))/1):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  m=1
        M15 N$98 VI- N$23 N$23 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        C7 N$124 VI- 0.25P
        M21 VB3 VB3 N$167 GROUND n_18_mm l=Lcf w={{({Wcf/(2*(k-1))}/1)}}
+  ad={eval((1/2-trunc(1/2)==0)?(({({Wcf/(2*(k-1))}/1)}*5.4e-07)/2):(({({Wcf/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wcf/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wcf/(2*(k-1))}/1)}*4.9e-07+(1-2)/2*({({Wcf/(2*(k-1))}/1)}*5.4e-07))/1):(({({Wcf/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wcf/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wcf/(2*(k-1))}/1)}+5.4e-07):((2*({({Wcf/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wcf/(2*(k-1))}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wcf/(2*(k-1))}/1)}+4.9e-07)+(1-2)*({({Wcf/(2*(k-1))}/1)}+5.4e-07))/1):((2*({({Wcf/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wcf/(2*(k-1))}/1)}+5.4e-07))/1))}
+  m=1
        M6 VO+ VB3 N$103 GROUND n_18_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*5.4e-07)/2):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*4.9e-07+(1-2)/2*({(Wcf/1)}*5.4e-07))/1):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+5.4e-07):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+4.9e-07)+(1-2)*({(Wcf/1)}+5.4e-07))/1):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  m=1
        M3A N$5 N$98 GROUND GROUND n_18_mm l=Lf w={{({k*Wf}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({k*Wf}/1)}*5.4e-07)/2):(({({k*Wf}/1)}*4.9e-07+((1-1)*{({k*Wf}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({k*Wf}/1)}*4.9e-07+(1-2)/2*({({k*Wf}/1)}*5.4e-07))/1):(({({k*Wf}/1)}*4.9e-07+((1-1)*{({k*Wf}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({k*Wf}/1)}+5.4e-07):((2*({({k*Wf}/1)}+4.9e-07)+(1-1)*({({k*Wf}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({k*Wf}/1)}+4.9e-07)+(1-2)*({({k*Wf}/1)}+5.4e-07))/1):((2*({({k*Wf}/1)}+4.9e-07)+(1-1)*({({k*Wf}/1)}+5.4e-07))/1))}
+  m=1
        M22 N$167 N$167 GROUND GROUND n_18_mm l={Lf} w={{({Wf/(2*(k-1))}/1)}}
+  ad={eval((1/2-trunc(1/2)==0)?(({({Wf/(2*(k-1))}/1)}*5.4e-07)/2):(({({Wf/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wf/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wf/(2*(k-1))}/1)}*4.9e-07+(1-2)/2*({({Wf/(2*(k-1))}/1)}*5.4e-07))/1):(({({Wf/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wf/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wf/(2*(k-1))}/1)}+5.4e-07):((2*({({Wf/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wf/(2*(k-1))}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wf/(2*(k-1))}/1)}+4.9e-07)+(1-2)*({({Wf/(2*(k-1))}/1)}+5.4e-07))/1):((2*({({Wf/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wf/(2*(k-1))}/1)}+5.4e-07))/1))}
+  m=1
        M3B N$47 N$98 GROUND GROUND n_18_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*5.4e-07)/2):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*4.9e-07+(1-2)/2*({(Wf/1)}*5.4e-07))/1):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+5.4e-07):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+4.9e-07)+(1-2)*({(Wf/1)}+5.4e-07))/1):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  m=1
        R4 VI- VO+ 100gig
        M7 VO- VB2 N$17 VDD p_18_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*5.4e-07)/2):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*4.9e-07+(1-2)/2*({(Wcl/1)}*5.4e-07))/1):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+5.4e-07):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+4.9e-07)+(1-2)*({(Wcl/1)}+5.4e-07))/1):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  m=1
        M16 N$103 VI- N$23 N$23 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M4 VB2 N$195 GROUND GROUND n_18_mm l=0.5u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        M1 VB3 VB1T VDD VDD p_18_mm l=0.5u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        V3 VDD GROUND DC 1.8V
        V2 VOCM GROUND DC 0.9
        R6 N$26 VI+ 100gig
        E5 N$42 N$41 Vo+ 0 0.5
        M18 N$103 N$105 GROUND GROUND n_18_mm l=Lf w={{({k*Wf}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({k*Wf}/1)}*5.4e-07)/2):(({({k*Wf}/1)}*4.9e-07+((1-1)*{({k*Wf}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({k*Wf}/1)}*4.9e-07+(1-2)/2*({({k*Wf}/1)}*5.4e-07))/1):(({({k*Wf}/1)}*4.9e-07+((1-1)*{({k*Wf}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({k*Wf}/1)}+5.4e-07):((2*({({k*Wf}/1)}+4.9e-07)+(1-1)*({({k*Wf}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({k*Wf}/1)}+4.9e-07)+(1-2)*({({k*Wf}/1)}+5.4e-07))/1):((2*({({k*Wf}/1)}+4.9e-07)+(1-1)*({({k*Wf}/1)}+5.4e-07))/1))}
+  m=1
        I1 VB1T GROUND DC Ib
        M25 VB2 VB2 N$181 VDD p_18_mm l=Lcl w={{({Wcl/(2*(k-1))}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wcl/(2*(k-1))}/1)}*5.4e-07)/2):(({({Wcl/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wcl/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wcl/(2*(k-1))}/1)}*4.9e-07+(1-2)/2*({({Wcl/(2*(k-1))}/1)}*5.4e-07))/1):(({({Wcl/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wcl/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wcl/(2*(k-1))}/1)}+5.4e-07):((2*({({Wcl/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wcl/(2*(k-1))}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wcl/(2*(k-1))}/1)}+4.9e-07)+(1-2)*({({Wcl/(2*(k-1))}/1)}+5.4e-07))/1):((2*({({Wcl/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wcl/(2*(k-1))}/1)}+5.4e-07))/1))}
+  m=1
        M26 N$181 N$181 VDD VDD p_18_mm l=Ll w={{({Wl/(2*(k-1))}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wl/(2*(k-1))}/1)}*5.4e-07)/2):(({({Wl/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wl/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wl/(2*(k-1))}/1)}*4.9e-07+(1-2)/2*({({Wl/(2*(k-1))}/1)}*5.4e-07))/1):(({({Wl/(2*(k-1))}/1)}*4.9e-07+((1-1)*{({Wl/(2*(k-1))}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wl/(2*(k-1))}/1)}+5.4e-07):((2*({({Wl/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wl/(2*(k-1))}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wl/(2*(k-1))}/1)}+4.9e-07)+(1-2)*({({Wl/(2*(k-1))}/1)}+5.4e-07))/1):((2*({({Wl/(2*(k-1))}/1)}+4.9e-07)+(1-1)*({({Wl/(2*(k-1))}/1)}+5.4e-07))/1))}
+  m=1
        M3 N$195 VB1T VDD VDD p_18_mm l=0.5u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        E7 VDD CMFB N$42 VOCM -30
        V1 N$29 GROUND PULSE ( -0.1V 0.1V 10nS 0.01nS 0.01nS 10nS 20nS )
        M0 N$23 VB1T VDD VDD p_18_mm l=0.5u w=64u ad=31.36p as=31.36p pd=0.129m
+  ps=0.129m m=1
        R5 N$124 VI- 100gig
        C6 VI- VO+ 1P
        M12 N$105 VB3 N$106 GROUND n_18_mm l=Laux w={{(Waux/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Waux/1)}*5.4e-07)/2):(({(Waux/1)}*4.9e-07+((1-1)*{(Waux/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Waux/1)}*4.9e-07+(1-2)/2*({(Waux/1)}*5.4e-07))/1):(({(Waux/1)}*4.9e-07+((1-1)*{(Waux/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Waux/1)}+5.4e-07):((2*({(Waux/1)}+4.9e-07)+(1-1)*({(Waux/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Waux/1)}+4.9e-07)+(1-2)*({(Waux/1)}+5.4e-07))/1):((2*({(Waux/1)}+4.9e-07)+(1-1)*({(Waux/1)}+5.4e-07))/1))}
+  m=1
        M17 N$106 N$105 GROUND GROUND n_18_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*5.4e-07)/2):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*4.9e-07+(1-2)/2*({(Wf/1)}*5.4e-07))/1):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+5.4e-07):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+4.9e-07)+(1-2)*({(Wf/1)}+5.4e-07))/1):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  m=1
        R3 VI+ VO- 100gig
        M1A N$5 VI+ N$23 N$23 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
*
.end
