*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Wed Oct 30 2013 at 15:21:04

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/OTA
*
        I3 VCASP VCASN DC Icas
        V4 VOCM GROUND DC 0.9
        C1 VI+ VI+ 0.1P
        M2 N$535 VI+ N$897 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M6 N$535 VB GROUND GROUND n_18_mm l=Llt w={{(Wlt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wlt/1)}*5.4e-07)/2):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wlt/1)}*4.9e-07+(1-2)/2*({(Wlt/1)}*5.4e-07))/1):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wlt/1)}+5.4e-07):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wlt/1)}+4.9e-07)+(1-2)*({(Wlt/1)}+5.4e-07))/1):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  m=1
        M11 VB VB GROUND GROUND n_18_mm l=Llt w={{(Wlt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wlt/1)}*5.4e-07)/2):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wlt/1)}*4.9e-07+(1-2)/2*({(Wlt/1)}*5.4e-07))/1):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wlt/1)}+5.4e-07):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wlt/1)}+4.9e-07)+(1-2)*({(Wlt/1)}+5.4e-07))/1):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  m=1
        M33 VO+ VCASN N$1070 GROUND n_18_mm l=Ll w={{(Wcasn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasn/1)}*5.4e-07)/2):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasn/1)}*4.9e-07+(1-2)/2*({(Wcasn/1)}*5.4e-07))/1):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasn/1)}+5.4e-07):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasn/1)}+4.9e-07)+(1-2)*({(Wcasn/1)}+5.4e-07))/1):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  m=1
        M5 N$536 VB GROUND GROUND n_18_mm l=Llt w={{(Wlt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wlt/1)}*5.4e-07)/2):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wlt/1)}*4.9e-07+(1-2)/2*({(Wlt/1)}*5.4e-07))/1):(({(Wlt/1)}*4.9e-07+((1-1)*{(Wlt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wlt/1)}+5.4e-07):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wlt/1)}+4.9e-07)+(1-2)*({(Wlt/1)}+5.4e-07))/1):((2*({(Wlt/1)}+4.9e-07)+(1-1)*({(Wlt/1)}+5.4e-07))/1))}
+  m=1
        M1 N$897 N$535 VDD VDD p_18_mm l=Lt w={{(Wt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wt/1)}*5.4e-07)/2):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wt/1)}*4.9e-07+(1-2)/2*({(Wt/1)}*5.4e-07))/1):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wt/1)}+5.4e-07):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wt/1)}+4.9e-07)+(1-2)*({(Wt/1)}+5.4e-07))/1):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  m=1
        M7 N$1239 VI+ N$654 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        V1 VDD GROUND DC 1.8V
        E5 GROUND CMFB N$821 VOCM 10
        M19 N$1242 CMFB GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        E3 N$830 GROUND Vo- 0 0.5
        C3 VOCM VO- 4P
        R3 VI- VI- 10gig
        R2 VI- VI- 10gig
        V2 N$1204 GROUND DC 0V AC 1 0
        C6 VI- VI- 0.1P
        M36 N$1078 N$1227 VDD VDD p_18_mm l=Loutp w={{({n*Wmp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({n*Wmp}/1)}*5.4e-07)/2):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({n*Wmp}/1)}*4.9e-07+(1-2)/2*({({n*Wmp}/1)}*5.4e-07))/1):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({n*Wmp}/1)}+5.4e-07):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({n*Wmp}/1)}+4.9e-07)+(1-2)*({({n*Wmp}/1)}+5.4e-07))/1):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  m=1
        M16 N$1242 N$1240 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M15 N$1120 VCASN GROUND GROUND n_18_mm l={{4*Ll}} w={{({k*Wl}/1)}}
+  ad={eval((1/2-trunc(1/2)==0)?(({({k*Wl}/1)}*5.4e-07)/2):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({k*Wl}/1)}*4.9e-07+(1-2)/2*({({k*Wl}/1)}*5.4e-07))/1):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({k*Wl}/1)}+5.4e-07):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({k*Wl}/1)}+4.9e-07)+(1-2)*({({k*Wl}/1)}+5.4e-07))/1):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  m=1
        I1 VDD VB DC Ib
        M3 N$654 N$536 VDD VDD p_18_mm l=Lt w={{(Wt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wt/1)}*5.4e-07)/2):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wt/1)}*4.9e-07+(1-2)/2*({(Wt/1)}*5.4e-07))/1):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wt/1)}+5.4e-07):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wt/1)}+4.9e-07)+(1-2)*({(Wt/1)}+5.4e-07))/1):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  m=1
        M9 N$1240 N$1223 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        E2 N$821 N$830 Vo+ 0 0.5
        M24 N$1242 N$1242 VDD VDD p_18_mm l=Loutp w={{(Wmp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wmp/1)}*5.4e-07)/2):(({(Wmp/1)}*4.9e-07+((1-1)*{(Wmp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wmp/1)}*4.9e-07+(1-2)/2*({(Wmp/1)}*5.4e-07))/1):(({(Wmp/1)}*4.9e-07+((1-1)*{(Wmp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wmp/1)}+5.4e-07):((2*({(Wmp/1)}+4.9e-07)+(1-1)*({(Wmp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wmp/1)}+4.9e-07)+(1-2)*({(Wmp/1)}+5.4e-07))/1):((2*({(Wmp/1)}+4.9e-07)+(1-1)*({(Wmp/1)}+5.4e-07))/1))}
+  m=1
        M13 VCASP VCASP N$1135 VDD p_18_mm l=Loutp w={{(Wcasp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasp/1)}*5.4e-07)/2):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasp/1)}*4.9e-07+(1-2)/2*({(Wcasp/1)}*5.4e-07))/1):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasp/1)}+5.4e-07):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasp/1)}+4.9e-07)+(1-2)*({(Wcasp/1)}+5.4e-07))/1):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  m=1
        V3 N$1249 GROUND PULSE ( -0.1V 0.1V 10nS 1nS 1nS 10nS 20nS )
        M35 VO- VCASP N$1078 VDD p_18_mm l=Loutp w={{(Wcasp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasp/1)}*5.4e-07)/2):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasp/1)}*4.9e-07+(1-2)/2*({(Wcasp/1)}*5.4e-07))/1):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasp/1)}+5.4e-07):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasp/1)}+4.9e-07)+(1-2)*({(Wcasp/1)}+5.4e-07))/1):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  m=1
        M17 N$1227 N$1239 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M31 N$1070 N$1239 GROUND GROUND n_18_mm l=Ll w={{({k*Wl}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({k*Wl}/1)}*5.4e-07)/2):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({k*Wl}/1)}*4.9e-07+(1-2)/2*({({k*Wl}/1)}*5.4e-07))/1):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({k*Wl}/1)}+5.4e-07):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({k*Wl}/1)}+4.9e-07)+(1-2)*({({k*Wl}/1)}+5.4e-07))/1):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  m=1
        M14 VCASN VCASN N$1120 GROUND n_18_mm l=Ll w={{(Wcasn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasn/1)}*5.4e-07)/2):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasn/1)}*4.9e-07+(1-2)/2*({(Wcasn/1)}*5.4e-07))/1):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasn/1)}+5.4e-07):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasn/1)}+4.9e-07)+(1-2)*({(Wcasn/1)}+5.4e-07))/1):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  m=1
        M32 VO- VCASN N$1069 GROUND n_18_mm l=Ll w={{(Wcasn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasn/1)}*5.4e-07)/2):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasn/1)}*4.9e-07+(1-2)/2*({(Wcasn/1)}*5.4e-07))/1):(({(Wcasn/1)}*4.9e-07+((1-1)*{(Wcasn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasn/1)}+5.4e-07):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasn/1)}+4.9e-07)+(1-2)*({(Wcasn/1)}+5.4e-07))/1):((2*({(Wcasn/1)}+4.9e-07)+(1-1)*({(Wcasn/1)}+5.4e-07))/1))}
+  m=1
        V6 N$1087 GROUND DC 0.9
        M34 VO+ VCASP N$1079 VDD p_18_mm l=Loutp w={{(Wcasp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcasp/1)}*5.4e-07)/2):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcasp/1)}*4.9e-07+(1-2)/2*({(Wcasp/1)}*5.4e-07))/1):(({(Wcasp/1)}*4.9e-07+((1-1)*{(Wcasp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcasp/1)}+5.4e-07):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcasp/1)}+4.9e-07)+(1-2)*({(Wcasp/1)}+5.4e-07))/1):((2*({(Wcasp/1)}+4.9e-07)+(1-1)*({(Wcasp/1)}+5.4e-07))/1))}
+  m=1
        X_S2D2 VI+ VI- N$1087 N$1204 GROUND S2D
        E4 VO GROUND VO- VO+ 1
        M30 N$1069 N$1240 GROUND GROUND n_18_mm l=Ll w={{({k*Wl}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({k*Wl}/1)}*5.4e-07)/2):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({k*Wl}/1)}*4.9e-07+(1-2)/2*({({k*Wl}/1)}*5.4e-07))/1):(({({k*Wl}/1)}*4.9e-07+((1-1)*{({k*Wl}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({k*Wl}/1)}+5.4e-07):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({k*Wl}/1)}+4.9e-07)+(1-2)*({({k*Wl}/1)}+5.4e-07))/1):((2*({({k*Wl}/1)}+4.9e-07)+(1-1)*({({k*Wl}/1)}+5.4e-07))/1))}
+  m=1
        M10 N$1239 N$1223 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M4 N$536 VI- N$654 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        R1 VI+ VI+ 10gig
        M12 N$1135 VCASP VDD VDD p_18_mm l={{4*Loutp}} w={{({n*Wmp}/1)}}
+  ad={eval((1/2-trunc(1/2)==0)?(({({n*Wmp}/1)}*5.4e-07)/2):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({n*Wmp}/1)}*4.9e-07+(1-2)/2*({({n*Wmp}/1)}*5.4e-07))/1):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({n*Wmp}/1)}+5.4e-07):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({n*Wmp}/1)}+4.9e-07)+(1-2)*({({n*Wmp}/1)}+5.4e-07))/1):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  m=1
        R4 VI+ VI+ 10gig
        M20 N$1227 CMFB GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M37 N$1079 N$1242 VDD VDD p_18_mm l=Loutp w={{({n*Wmp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({n*Wmp}/1)}*5.4e-07)/2):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({n*Wmp}/1)}*4.9e-07+(1-2)/2*({({n*Wmp}/1)}*5.4e-07))/1):(({({n*Wmp}/1)}*4.9e-07+((1-1)*{({n*Wmp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({n*Wmp}/1)}+5.4e-07):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({n*Wmp}/1)}+4.9e-07)+(1-2)*({({n*Wmp}/1)}+5.4e-07))/1):((2*({({n*Wmp}/1)}+4.9e-07)+(1-1)*({({n*Wmp}/1)}+5.4e-07))/1))}
+  m=1
        C4 VO+ VOCM 4P
        M8 N$1240 VI- N$897 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        C5 VI- VI- 0.1P
        C2 VI+ VI+ 0.1P
        R6 N$1223 N$1240 Rr
        R5 N$1239 N$1223 Rr
        M25 N$1227 N$1227 VDD VDD p_18_mm l=Loutp w={{(Wmp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wmp/1)}*5.4e-07)/2):(({(Wmp/1)}*4.9e-07+((1-1)*{(Wmp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wmp/1)}*4.9e-07+(1-2)/2*({(Wmp/1)}*5.4e-07))/1):(({(Wmp/1)}*4.9e-07+((1-1)*{(Wmp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wmp/1)}+5.4e-07):((2*({(Wmp/1)}+4.9e-07)+(1-1)*({(Wmp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wmp/1)}+4.9e-07)+(1-2)*({(Wmp/1)}+5.4e-07))/1):((2*({(Wmp/1)}+4.9e-07)+(1-1)*({(Wmp/1)}+5.4e-07))/1))}
+  m=1
*
.end
