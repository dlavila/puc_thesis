*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Tue Nov  5 2013 at 10:30:35

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/folded_180
*
        C1 VI+ N$142 1P
        M14 VB3 VB3 VB4 GROUND n_18_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*5.4e-07)/2):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*4.9e-07+(1-2)/2*({(Wcf/1)}*5.4e-07))/1):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+5.4e-07):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+4.9e-07)+(1-2)*({(Wcf/1)}+5.4e-07))/1):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  m=1
        M9 VB4 VB4 GROUND GROUND n_18_mm l=Lf w={{({Wf/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wf/2}/1)}*5.4e-07)/2):(({({Wf/2}/1)}*4.9e-07+((1-1)*{({Wf/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wf/2}/1)}*4.9e-07+(1-2)/2*({({Wf/2}/1)}*5.4e-07))/1):(({({Wf/2}/1)}*4.9e-07+((1-1)*{({Wf/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wf/2}/1)}+5.4e-07):((2*({({Wf/2}/1)}+4.9e-07)+(1-1)*({({Wf/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wf/2}/1)}+4.9e-07)+(1-2)*({({Wf/2}/1)}+5.4e-07))/1):((2*({({Wf/2}/1)}+4.9e-07)+(1-1)*({({Wf/2}/1)}+5.4e-07))/1))}
+  m=1
        I4 VB2 VB3 DC 35u
        V4 N$28 GROUND DC 0V AC 1 0
        M11 N$137 VB4 GROUND GROUND n_18_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*5.4e-07)/2):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*4.9e-07+(1-2)/2*({(Wf/1)}*5.4e-07))/1):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+5.4e-07):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+4.9e-07)+(1-2)*({(Wf/1)}+5.4e-07))/1):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  m=1
        M10 N$124 VB1T VDD VDD p_18_mm l=1u w=100u ad=49p as=49p pd=0.201m
+  ps=0.201m m=1
        C5 VI- N$153 1P
        M12 N$131 VI+ N$124 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M13 VB1T VB1T VDD VDD p_18_mm l=1u w=14u ad=6.86p as=6.86p pd=28.98u
+  ps=28.98u m=1
        I2 VB1T GROUND DC 10u
        E5 VDD CMFB N$39 VOCM -10
        E3 N$38 GROUND Vo- 0 0.5
        E2 N$39 N$38 Vo+ 0 0.5
        C4 VO+ VOCM 4P
        C3 VOCM VO- 4P
        V2 VOCM GROUND DC 0.9
        R4 VI+ VI+ 100gig
        R3 VI- VI- 100gig
        R2 VI- N$153 100gig
        R1 VI+ N$142 100gig
        C7 VI- VI- 0.25P
        M15 VB2 VB2 N$141 VDD p_18_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*5.4e-07)/2):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*4.9e-07+(1-2)/2*({(Wcl/1)}*5.4e-07))/1):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+5.4e-07):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+4.9e-07)+(1-2)*({(Wcl/1)}+5.4e-07))/1):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  m=1
        M16 N$141 N$141 VDD VDD p_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M7 VO- VB3 N$131 GROUND n_18_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*5.4e-07)/2):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*4.9e-07+(1-2)/2*({(Wcf/1)}*5.4e-07))/1):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+5.4e-07):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+4.9e-07)+(1-2)*({(Wcf/1)}+5.4e-07))/1):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  m=1
        V6 N$27 GROUND DC 0.9
        X_S2D2 VI+ VI- N$27 N$28 GROUND S2D
        C2 VI+ VI+ 0.25P
        M8 VO+ VB3 N$137 GROUND n_18_mm l=Lcf w={{(Wcf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcf/1)}*5.4e-07)/2):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcf/1)}*4.9e-07+(1-2)/2*({(Wcf/1)}*5.4e-07))/1):(({(Wcf/1)}*4.9e-07+((1-1)*{(Wcf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcf/1)}+5.4e-07):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcf/1)}+4.9e-07)+(1-2)*({(Wcf/1)}+5.4e-07))/1):((2*({(Wcf/1)}+4.9e-07)+(1-1)*({(Wcf/1)}+5.4e-07))/1))}
+  m=1
        E4 VO GROUND VO- VO+ 1
        M4 VO+ VB2 N$130 VDD p_18_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*5.4e-07)/2):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*4.9e-07+(1-2)/2*({(Wcl/1)}*5.4e-07))/1):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+5.4e-07):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+4.9e-07)+(1-2)*({(Wcl/1)}+5.4e-07))/1):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  m=1
        M3 N$130 CMFB VDD VDD p_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M1 N$137 VI- N$124 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M5 VO- VB2 N$128 VDD p_18_mm l=Lcl w={{(Wcl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wcl/1)}*5.4e-07)/2):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wcl/1)}*4.9e-07+(1-2)/2*({(Wcl/1)}*5.4e-07))/1):(({(Wcl/1)}*4.9e-07+((1-1)*{(Wcl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wcl/1)}+5.4e-07):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wcl/1)}+4.9e-07)+(1-2)*({(Wcl/1)}+5.4e-07))/1):((2*({(Wcl/1)}+4.9e-07)+(1-1)*({(Wcl/1)}+5.4e-07))/1))}
+  m=1
        M2 N$128 CMFB VDD VDD p_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        V3 VDD GROUND DC 1.8V
        M6 N$131 VB4 GROUND GROUND n_18_mm l=Lf w={{(Wf/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wf/1)}*5.4e-07)/2):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wf/1)}*4.9e-07+(1-2)/2*({(Wf/1)}*5.4e-07))/1):(({(Wf/1)}*4.9e-07+((1-1)*{(Wf/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wf/1)}+5.4e-07):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wf/1)}+4.9e-07)+(1-2)*({(Wf/1)}+5.4e-07))/1):((2*({(Wf/1)}+4.9e-07)+(1-1)*({(Wf/1)}+5.4e-07))/1))}
+  m=1
*
.end
