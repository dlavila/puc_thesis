*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Mon Jan 13 2014 at 17:18:30

*
* Globals.
*
.global VDD GROUND


*
* Component pathname : $MGC_DESIGN_KIT/symbols/MIMCAPS_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/MIMCAPS_MM/mimcaps_mm


*
* Component pathname : $MGC_DESIGN_KIT/symbols/RNHR1000_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/RNHR1000_MM/rnhr1000_mm

*
* Component pathname : $UTILS/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $SC_filter/default.group/logic.views/BUFFER
*
.subckt BUFFER  VO AGND AVDD VB1 VB2 VB3 VB4 VI+ VI- VNCAS VPCAS

        XR1 ND9 N$941 AVDD rnhr1000_mm lr=10u wr=2u m=1
        M64 ND1 N$752 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M14 ND7 VPCAS ND9 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M18 ND3 VI- N$209 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.744p
+  pd=3.04u ps=3.408u m=16
        M5 ND1 ND8 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p pd=3.04u
+  ps=4.51u m=4
        M8 ND8 VNCAS ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M2 N$165 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p
+  pd=2.14u ps=3.16u m=4
        M41 ND4 VI+ N$209 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.744p
+  pd=3.04u ps=3.408u m=16
        M42 N$427 N$427 N$209 AVDD p_18_mm l=0.45u w=8u ad=2.16p as=2.512p
+  pd=8.54u ps=10.228u m=10
        MOUTP VO ND9 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.702p
+  pd=3.04u ps=3.187u m=40
        M52 ND1 N$749 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        MIN1 ND1 VI- N$204 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.52p
+  pd=2.14u ps=2.65u m=8
        M1 N$209 VB2 N$206 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M11 ND9 VNCAS ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M9 ND6 VB3 ND3 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p pd=2.14u
+  ps=3.16u m=4
        M16 ND4 ND6 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        MOUTN VO ND7 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.467p
+  pd=2.14u ps=2.344u m=20
        M79 ND8 N$761 ND8 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M81 ND6 N$768 ND6 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M78 ND7 N$758 ND7 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M77 ND6 N$755 ND6 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M4 N$204 VB3 N$165 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p
+  pd=2.14u ps=3.16u m=4
        M10 ND8 VB2 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M80 ND9 N$764 ND9 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M90 ND7 N$801 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        XC1 N$943 VO mimcaps_mm w=13u l=6.5u m=6
        M51 ND1 N$688 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        XR4 ND7 N$943 AVDD rnhr1000_mm lr=10u wr=2u m=1
        XR3 ND7 N$943 AVDD rnhr1000_mm lr=10u wr=2u m=1
        XR2 ND9 N$941 AVDD rnhr1000_mm lr=10u wr=2u m=1
        M15 ND3 ND6 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        M13 ND6 VPCAS ND8 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M7 ND7 VB3 ND4 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.608p pd=2.14u
+  ps=3.16u m=4
        M67 ND8 N$812 ND8 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M68 ND9 N$816 ND9 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M12 ND9 VB2 ND2 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M50 N$427 N$427 N$204 AGND n_18_mm l=0.45u w=5.12u ad=1.382p as=1.608p
+  pd=5.66u ps=6.772u m=10
        M89 ND6 N$798 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M88 ND7 N$795 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M87 ND6 N$792 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M86 ND7 N$789 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M84 ND6 N$786 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M85 ND7 N$780 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M83 ND6 N$774 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M19 N$427 N$427 N$209 AVDD p_18_mm l=0.45u w=8u ad=2.16p as=2.512p
+  pd=8.54u ps=10.228u m=10
        XC2 N$941 VO mimcaps_mm w=13u l=6.5u m=6
        M66 ND7 N$702 ND7 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M65 ND6 N$672 ND6 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M63 ND1 N$668 ND1 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M3 N$206 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.812p
+  pd=3.04u ps=3.775u m=8
        M17 ND2 VI+ N$204 AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.52p
+  pd=2.14u ps=2.65u m=8
        M6 ND2 ND8 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p pd=3.04u
+  ps=4.51u m=4
        M55 ND8 N$695 ND8 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M56 ND9 N$650 ND9 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M82 ND7 N$771 ND7 AVDD p_18_mm l=0.45u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
.ends BUFFER

*
* Component pathname : $SC_filter/default.group/logic.views/BIAS_BUFFER
*
.subckt BIAS_BUFFER  VB1 VB2 VB3 VB4 VNCAS VPCAS AGND AVDD IB

        M74 VB3 N$65 VB3 AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M73 VB3 N$63 VB3 AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M48 IB IB AVDD AVDD p_18_mm l=0.45u w=5u ad=2.45p as=2.45p pd=10.98u
+  ps=10.98u m=1
        M45 VB3 IB AVDD AVDD p_18_mm l=0.45u w=5u ad=1.35p as=1.9p pd=5.54u
+  ps=8.26u m=4
        M43 VB4 IB AVDD AVDD p_18_mm l=0.45u w=5u ad=1.35p as=1.9p pd=5.54u
+  ps=8.26u m=4
        M22 VB2 VB2 N$54 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M40 VB1 VB2 N$60 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M38 N$60 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M37 N$59 VB1 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M39 VNCAS VB2 N$59 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M32 VNCAS VNCAS N$52 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M31 N$58 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M30 VB1 VB3 N$58 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M29 N$57 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M28 VB2 VB3 N$57 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M27 N$56 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M26 VPCAS VB3 N$56 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M25 N$55 VB4 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M36 N$54 VB2 AVDD AVDD p_18_mm l=2.25u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
        M24 N$53 VB3 AGND AGND n_18_mm l=2.25u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M21 VB3 VB3 N$53 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M35 N$52 N$52 AGND AGND n_18_mm l=0.45u w=1.6u ad=0.432p as=0.784p
+  pd=2.14u ps=4.18u m=2
        M23 VB4 VB3 N$55 AGND n_18_mm l=0.45u w=1.6u ad=0.784p as=0.784p
+  pd=4.18u ps=4.18u m=1
        M34 N$51 N$51 AVDD AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=0.95p
+  pd=3.04u ps=4.51u m=4
        M33 VPCAS VPCAS N$51 AVDD p_18_mm l=0.45u w=2.5u ad=0.675p as=1.225p
+  pd=3.04u ps=5.98u m=2
.ends BIAS_BUFFER

*
* MAIN CELL: Component pathname : $SC_filter/default.group/logic.views/testBuffer
*
        X_S2D1 N$46 N$78 N$29 N$31 GROUND S2D
        X_BUFFER1 VO GROUND VDD N$65 N$64 N$63 N$62 N$46 N$78 N$61 N$60 BUFFER
        X_BIAS_BUFFER1 N$65 N$64 N$63 N$62 N$61 N$60 GROUND VDD N$2 BIAS_BUFFER
        V3 N$31 GROUND DC 0V AC 1 0
        V2 N$29 GROUND DC 0.9V
        C1 VO GROUND 4P
        V1 VDD GROUND DC 1.8V
        I1 N$2 GROUND DC 3.75uA
*
.end
