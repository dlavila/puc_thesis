*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Tue Nov  5 2013 at 19:06:15

*
* Globals.
*
.global GROUND

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/noise_test
*
        M1 N$6 VI GROUND GROUND n_18_mm l=0.18u w=50u ad=24.5p as=24.5p
+  pd=0.101m ps=0.101m m=1
        H1 VO GROUND V2 -1
        V3 N$12 GROUND DC 0.7V
        V1 VI N$12 DC 0V AC 1 0
        V2 N$6 GROUND DC 1.8V
*
.end
