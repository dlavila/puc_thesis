*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Wed Dec 18 2013 at 14:58:36

*
* Globals.
*
.global VDD LS_BUFFER_VDD GROUND

*
* Component pathname : $SC_filter/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $LS_BUFFER/default.group/logic.views/LS_BUFFER_switch_X4
*
.subckt LS_BUFFER_SWITCH_X4  OUT E IN

        M12 OUT N$40 IN LS_BUFFER_VDD p_18_mm l=0.18u w=1.5u ad=0.405p as=0.488p
+  pd=2.04u ps=2.525u m=8
        M11 OUT E IN GROUND n_18_mm l=0.18u w=0.5u ad=0.135p as=0.163p pd=1.04u
+  ps=1.275u m=8
        M2 N$40 E LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=1.5u ad=0.405p
+  as=0.735p pd=2.04u ps=3.98u m=2
        M1 N$40 E GROUND GROUND n_18_mm l=0.18u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
.ends LS_BUFFER_SWITCH_X4

*
* Component pathname : $LS_BUFFER/default.group/logic.views/LS_BUFFER_inv_X4
*
.subckt LS_BUFFER_INV_X4  O I

        M2 O I LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=0.75u ad=0.203p
+  as=0.285p pd=1.29u ps=1.885u m=4
        M1 O I GROUND GROUND n_18_mm l=0.18u w=0.25u ad=67.5f as=95f pd=0.79u
+  ps=1.135u m=4
.ends LS_BUFFER_INV_X4

*
* Component pathname : $LS_BUFFER/default.group/logic.views/PHASE_GEN_nand_X4
*
.subckt PHASE_GEN_NAND_X4  O A B

        M1 O B LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=0.75u ad=0.203p
+  as=0.285p pd=1.29u ps=1.885u m=4
        M4 O A LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=0.75u ad=0.203p
+  as=0.285p pd=1.29u ps=1.885u m=4
        M3 N$75 B GROUND GROUND n_18_mm l=0.18u w=0.25u ad=67.5f as=95f
+  pd=0.79u ps=1.135u m=4
        M2 O A N$75 GROUND n_18_mm l=0.18u w=0.25u ad=67.5f as=95f pd=0.79u
+  ps=1.135u m=4
.ends PHASE_GEN_NAND_X4

*
* Component pathname : $LS_BUFFER/default.group/logic.views/LS_BUFFER_inv_X2
*
.subckt LS_BUFFER_INV_X2  O I

        M2 O I LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=0.75u ad=0.203p
+  as=0.368p pd=1.29u ps=2.48u m=2
        M1 O I GROUND GROUND n_18_mm l=0.18u w=0.25u ad=67.5f as=0.122p
+  pd=0.79u ps=1.48u m=2
.ends LS_BUFFER_INV_X2

*
* Component pathname : $LS_BUFFER/default.group/logic.views/PHASE_GEN
*
.subckt PHASE_GEN  PHI1 PHI2 CLK

        X_LS_BUFFER_INV_X46 PHI2 N$226 LS_BUFFER_INV_X4
        X_LS_BUFFER_INV_X45 N$226 N$225 LS_BUFFER_INV_X4
        X_LS_BUFFER_INV_X41 N$225 N$224 LS_BUFFER_INV_X4
        X_LS_BUFFER_INV_X44 PHI1 N$223 LS_BUFFER_INV_X4
        X_LS_BUFFER_INV_X42 N$221 N$9 LS_BUFFER_INV_X4
        X_LS_BUFFER_INV_X43 N$223 N$221 LS_BUFFER_INV_X4
        X_PHASE_GEN_NAND_X42 N$224 N$220 N$223 PHASE_GEN_NAND_X4
        X_LS_BUFFER_INV_X21 N$220 CLK LS_BUFFER_INV_X2
        X_PHASE_GEN_NAND_X41 N$9 CLK N$226 PHASE_GEN_NAND_X4
.ends PHASE_GEN

*
* Component pathname : $LS_BUFFER/default.group/logic.views/LS_BUFFER_inv_X8
*
.subckt LS_BUFFER_INV_X8  O I

        M2 O I LS_BUFFER_VDD LS_BUFFER_VDD p_18_mm l=0.18u w=0.75u ad=0.203p
+  as=0.244p pd=1.29u ps=1.588u m=8
        M1 O I GROUND GROUND n_18_mm l=0.18u w=0.25u ad=67.5f as=81.25f
+  pd=0.79u ps=0.963u m=8
.ends LS_BUFFER_INV_X8

*
* MAIN CELL: Component pathname : $LS_BUFFER/default.group/logic.views/LS_BUFFER
*
        V6 N$878 GROUND DC 0.9V
        X_S2D1 V+ V- N$878 VI GROUND S2D
        V9 N$938 GROUND DC 1V
        I2 N$985 GROUND DC Ib
        M17 N$983 N$983 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        X_LS_BUFFER_SWITCH_X41 V+ PHI1 N$921 LS_BUFFER_SWITCH_X4
        M24 N$988 N$994 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M23 VO+ N$993 VDD VDD p_18_mm l=Lp w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M15 N$978 N$984 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M16 N$984 N$984 GROUND GROUND n_18_mm l=Ln w={{({Wn/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/5}/1)}*5.4e-07)/2):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/5}/1)}*4.9e-07+(1-2)/2*({({Wn/5}/1)}*5.4e-07))/1):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/5}/1)}+5.4e-07):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/5}/1)}+4.9e-07)+(1-2)*({({Wn/5}/1)}+5.4e-07))/1):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  m=1
        E1 VI+ GROUND N$924 GROUND 1
        X_PHASE_GEN1 N$951 N$952 N$207 PHASE_GEN
        X_LS_BUFFER_SWITCH_X46 N$936 PHI2 N$938 LS_BUFFER_SWITCH_X4
        V5 N$207 GROUND PULSE ( 0V 1.8V 10nS 0.1nS 0.1nS 10nS 20nS )
        M18 N$985 N$985 N$983 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M14 VO- N$983 VDD VDD p_18_mm l=Lp w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M29 N$994 N$995 N$996 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M28 N$996 N$993 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        E4 VI_I GROUND VI+ VI- 1
        V3 VDD GROUND DC 1.8V
        M13 VO- N$978 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M12 N$978 VI- VO- VO- p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        V8 N$242 GROUND DC 1V
        E2 VO GROUND VO+ VO- 1
        C1 N$921 N$924 4.9P
        V1 N$920 N$242 DC -0.1V
        E3 VI- GROUND N$936 GROUND 1
        V2 VI GROUND SIN ( 0 0.1v 5Meg 0 0 )
        X_LS_BUFFER_SWITCH_X44 V- PHI1 N$940 LS_BUFFER_SWITCH_X4
        C4 N$940 N$936 4.9P
        V7 N$942 N$938 DC -0.1V
        M27 N$995 N$995 N$993 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        I3 N$995 GROUND DC Ib
        M26 N$993 N$993 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M25 N$994 N$994 GROUND GROUND n_18_mm l=Ln w={{({Wn/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/5}/1)}*5.4e-07)/2):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/5}/1)}*4.9e-07+(1-2)/2*({({Wn/5}/1)}*5.4e-07))/1):(({({Wn/5}/1)}*4.9e-07+((1-1)*{({Wn/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/5}/1)}+5.4e-07):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/5}/1)}+4.9e-07)+(1-2)*({({Wn/5}/1)}+5.4e-07))/1):((2*({({Wn/5}/1)}+4.9e-07)+(1-1)*({({Wn/5}/1)}+5.4e-07))/1))}
+  m=1
        X_LS_BUFFER_INV_X84 PHI1 N$960 LS_BUFFER_INV_X8
        X_LS_BUFFER_INV_X83 N$960 N$952 LS_BUFFER_INV_X8
        X_LS_BUFFER_INV_X82 PHI2 N$959 LS_BUFFER_INV_X8
        X_LS_BUFFER_INV_X81 N$959 N$951 LS_BUFFER_INV_X8
        M22 VO+ N$988 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M21 N$988 VI+ VO+ VO+ p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M20 N$984 N$985 N$986 VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        M19 N$986 N$983 VDD VDD p_18_mm l=Lp w={{({Wp/5}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/5}/1)}*5.4e-07)/2):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/5}/1)}*4.9e-07+(1-2)/2*({({Wp/5}/1)}*5.4e-07))/1):(({({Wp/5}/1)}*4.9e-07+((1-1)*{({Wp/5}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/5}/1)}+5.4e-07):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/5}/1)}+4.9e-07)+(1-2)*({({Wp/5}/1)}+5.4e-07))/1):((2*({({Wp/5}/1)}+4.9e-07)+(1-1)*({({Wp/5}/1)}+5.4e-07))/1))}
+  m=1
        X_LS_BUFFER_SWITCH_X45 N$940 PHI2 N$942 LS_BUFFER_SWITCH_X4
        X_LS_BUFFER_SWITCH_X43 N$924 PHI2 N$242 LS_BUFFER_SWITCH_X4
        X_LS_BUFFER_SWITCH_X42 N$921 PHI2 N$920 LS_BUFFER_SWITCH_X4
        V4 LS_BUFFER_VDD GROUND DC 1.8V
*
.end
