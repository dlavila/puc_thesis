*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Fri Oct 25 2013 at 17:30:14

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/OTA2
*
        M8 VO2 N$71 VDD VDD p_18_mm l=Lin w={{({4*Win}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({4*Win}/1)}*5.4e-07)/2):(({({4*Win}/1)}*4.9e-07+((1-1)*{({4*Win}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({4*Win}/1)}*4.9e-07+(1-2)/2*({({4*Win}/1)}*5.4e-07))/1):(({({4*Win}/1)}*4.9e-07+((1-1)*{({4*Win}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({4*Win}/1)}+5.4e-07):((2*({({4*Win}/1)}+4.9e-07)+(1-1)*({({4*Win}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({4*Win}/1)}+4.9e-07)+(1-2)*({({4*Win}/1)}+5.4e-07))/1):((2*({({4*Win}/1)}+4.9e-07)+(1-1)*({({4*Win}/1)}+5.4e-07))/1))}
+  m=1
        M7 VO2 VO GROUND GROUND n_18_mm l=Ll w={{({4*Wl}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({4*Wl}/1)}*5.4e-07)/2):(({({4*Wl}/1)}*4.9e-07+((1-1)*{({4*Wl}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({4*Wl}/1)}*4.9e-07+(1-2)/2*({({4*Wl}/1)}*5.4e-07))/1):(({({4*Wl}/1)}*4.9e-07+((1-1)*{({4*Wl}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({4*Wl}/1)}+5.4e-07):((2*({({4*Wl}/1)}+4.9e-07)+(1-1)*({({4*Wl}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({4*Wl}/1)}+4.9e-07)+(1-2)*({({4*Wl}/1)}+5.4e-07))/1):((2*({({4*Wl}/1)}+4.9e-07)+(1-1)*({({4*Wl}/1)}+5.4e-07))/1))}
+  m=1
        M6 N$71 N$71 VDD VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M5 N$22 N$71 VDD VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M2 N$47 N$47 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        M1 VO N$47 GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        V2 N$27 GROUND DC Vicm
        X_S2D1 VI+ VI- N$27 N$28 GROUND S2D
        V1 VDD GROUND DC 1.8V
        V3 N$28 GROUND DC 0V AC 1 0
        I1 N$71 GROUND DC 100u
        M3 VO VI- N$22 N$22 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M4 N$47 VI+ N$22 N$22 p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
*
.end
