*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Wed Oct 30 2013 at 18:03:55

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCN_Bias
*
.subckt AUX_FCN_BIAS  VB1 VB2 VB3 VB4 IIN VDD VSS

        M7 N$15 VB1 VDD VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M6 VB1 VB2 N$15 VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M5 VB2 VB2 N$14 VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M3 N$14 VB2 VDD VDD p_18_mm l=2.5u w=0.24u ad=0.118p as=0.118p pd=1.46u
+  ps=1.46u m=1
        M22 N$16 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M12 N$13 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M11 VB4 VB3 N$13 VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M9 N$12 VB3 VSS VSS n_18_mm l=2.5u w=0.75u ad=0.368p as=0.368p pd=2.48u
+  ps=2.48u m=1
        M8 VB3 VB3 N$12 VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M18 VB4 IIN N$11 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M16 N$11 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M25 N$10 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M24 VB3 IIN N$10 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M27 N$17 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M29 N$8 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p pd=3.38u
+  ps=3.38u m=1
        M28 IIN IIN N$8 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p pd=3.38u
+  ps=3.38u m=1
        M26 VB1 VB3 N$17 VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M23 VB2 VB3 N$16 VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
.ends AUX_FCN_BIAS

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCN
*
.subckt AUX_FCN  VO VB1 VB2 VB3 VB4 VDD VI+ VI- VSS

        M19 N$681 VB1 VDD VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M10 VO VB3 N$614 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M20 N$616 N$678 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M21 N$678 VB3 N$616 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M2 N$677 VI+ N$619 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M15 VO VB2 N$681 VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M17 N$614 N$678 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M13 N$677 VB1 VDD VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M4 N$619 VB4 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M1 N$681 VI- N$619 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M14 N$678 VB2 N$677 VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
.ends AUX_FCN

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCP
*
.subckt AUX_FCP  VO VB1 VB2 VB3 VB4 VDD VI+ VI- VSS

        M6 N$252 VB1 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M15 VO VB2 N$248 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M14 N$249 VB2 N$246 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M13 N$246 N$249 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M19 N$248 N$249 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M30 N$251 VI- N$252 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M20 VO VB3 N$251 VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M21 N$251 VB4 VSS VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M17 N$249 VB3 N$253 VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M3 N$253 VI+ N$252 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M10 N$253 VB4 VSS VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
.ends AUX_FCP

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCP_Bias
*
.subckt AUX_FCP_BIAS  VB1 VB2 VB3 VB4 IIN VDD VSS

        M12 VB1 VB3 N$32 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M7 N$32 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M4 N$31 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M2 VB2 VB3 N$31 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M1 VB2 VB2 N$33 VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M11 N$30 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M8 VB4 VB3 N$30 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M5 N$29 VB3 VSS VSS n_18_mm l=2.5u w=0.24u ad=0.118p as=0.118p pd=1.46u
+  ps=1.46u m=1
        M9 VB3 VB3 N$29 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M18 VB4 IIN N$25 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M16 N$25 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M25 N$24 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M24 VB3 IIN N$24 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M23 N$34 VB1 VDD VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M29 N$22 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M28 IIN IIN N$22 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M26 VB1 VB2 N$34 VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M22 N$33 VB2 VDD VDD p_18_mm l=2.5u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
.ends AUX_FCP_BIAS

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/Tel_OTA
*
        R3 N$419 VI- 10gig
        V2 VDD GROUND DC 1.8V
        R6 VOCM VDD 10gig
        M28 N$782 N$782 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M26 N$781 N$781 N$782 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        I1 N$781 VB4 DC Ib
        I2 IREFN GROUND DC Iref
        M2 VO- N$774 N$775 N$776 n_18_mm l=Ln w={{(Wncas/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wncas/1)}*5.4e-07)/2):(({(Wncas/1)}*4.9e-07+((1-1)*{(Wncas/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wncas/1)}*4.9e-07+(1-2)/2*({(Wncas/1)}*5.4e-07))/1):(({(Wncas/1)}*4.9e-07+((1-1)*{(Wncas/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wncas/1)}+5.4e-07):((2*({(Wncas/1)}+4.9e-07)+(1-1)*({(Wncas/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wncas/1)}+4.9e-07)+(1-2)*({(Wncas/1)}+5.4e-07))/1):((2*({(Wncas/1)}+4.9e-07)+(1-1)*({(Wncas/1)}+5.4e-07))/1))}
+  m=1
        M44 N$794 N$785 N$793 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M43 N$793 N$788 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M42 VCASP N$791 VDD VDD p_18_mm l=2.2u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M41 N$791 N$791 VCASP VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M39 N$791 N$785 N$790 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M5 N$779 VI- N$776 N$776 n_18_mm l=0.18u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        X_AUX_FCN_BIAS1 N$83 N$93 N$94 N$95 IREFN VDD GROUND AUX_FCN_BIAS
        M34 VCASN N$785 GROUND GROUND n_18_mm l=2.2u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        V1 N$767 GROUND DC 0V AC 1 0
        X_AUX_FCN2 N$762 N$83 N$93 N$94 N$95 VDD VCASP N$725 GROUND AUX_FCN
        C6 N$419 VI- 0.1P
        C5 VI- VO+ 0.1P
        M47 VB4 VB4 GROUND GROUND n_18_mm l=0.45u w={{({Wn/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/2}/1)}*5.4e-07)/2):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/2}/1)}*4.9e-07+(1-2)/2*({({Wn/2}/1)}*5.4e-07))/1):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/2}/1)}+5.4e-07):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/2}/1)}+4.9e-07)+(1-2)*({({Wn/2}/1)}+5.4e-07))/1):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  m=1
        M46 N$795 N$794 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M45 N$794 N$791 N$795 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        X_AUX_FCP1 N$778 N$64 N$63 N$62 N$61 VDD VCASN N$779 GROUND AUX_FCP
        X_S2D2 N$633 N$419 VOCM N$754 GROUND S2D
        E5 VDD CMFB N$187 VOCM -30
        C1 N$633 VI+ 0.1P
        M9 N$725 CMFB VDD VDD p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        C2 VI+ VO- 0.1P
        X_AUX_FCN1 N$764 N$83 N$93 N$94 N$95 VDD VCASP N$716 GROUND AUX_FCN
        M38 N$790 N$788 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M37 N$789 N$788 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M36 N$788 N$785 N$789 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M3 VO- N$762 N$725 VDD p_18_mm l=Lp w={{(Wpcas/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wpcas/1)}*5.4e-07)/2):(({(Wpcas/1)}*4.9e-07+((1-1)*{(Wpcas/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wpcas/1)}*4.9e-07+(1-2)/2*({(Wpcas/1)}*5.4e-07))/1):(({(Wpcas/1)}*4.9e-07+((1-1)*{(Wpcas/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wpcas/1)}+5.4e-07):((2*({(Wpcas/1)}+4.9e-07)+(1-1)*({(Wpcas/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wpcas/1)}+4.9e-07)+(1-2)*({(Wpcas/1)}+5.4e-07))/1):((2*({(Wpcas/1)}+4.9e-07)+(1-1)*({(Wpcas/1)}+5.4e-07))/1))}
+  m=1
        M6 N$776 VB4 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        R1 VI+ VO- 10gig
        C10 N$764 VDD Cc
        C9 GROUND N$778 Cc
        C8 N$762 VDD Cc
        C7 GROUND N$774 Cc
        E3 N$188 GROUND Vo- 0 0.5
        C4 VO+ VOCM 0.1P
        I3 IREFP GROUND DC Iref
        R5 GROUND VOCM 10gig
        X_AUX_FCP2 N$774 N$64 N$63 N$62 N$61 VDD VCASN N$775 GROUND AUX_FCP
        V7 N$754 GROUND PULSE ( -0.5V 0.5V 10nS 0.01nS 0.01nS 10nS 20nS
+  )
        E2 N$187 N$188 Vo+ 0 0.5
        X_AUX_FCP_BIAS1 N$64 N$63 N$62 N$61 IREFP VDD GROUND AUX_FCP_BIAS
        C3 VOCM VO- 0.1P
        M8 N$716 CMFB VDD VDD p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        R2 VI- VO+ 10gig
        R4 N$633 VI+ 10gig
        M33 N$788 N$781 N$786 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M32 N$786 N$782 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M31 N$785 N$785 VCASN GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M30 N$783 N$782 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M29 N$785 N$781 N$783 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M4 VO+ N$764 N$716 VDD p_18_mm l=Lp w={{(Wpcas/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wpcas/1)}*5.4e-07)/2):(({(Wpcas/1)}*4.9e-07+((1-1)*{(Wpcas/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wpcas/1)}*4.9e-07+(1-2)/2*({(Wpcas/1)}*5.4e-07))/1):(({(Wpcas/1)}*4.9e-07+((1-1)*{(Wpcas/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wpcas/1)}+5.4e-07):((2*({(Wpcas/1)}+4.9e-07)+(1-1)*({(Wpcas/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wpcas/1)}+4.9e-07)+(1-2)*({(Wpcas/1)}+5.4e-07))/1):((2*({(Wpcas/1)}+4.9e-07)+(1-1)*({(Wpcas/1)}+5.4e-07))/1))}
+  m=1
        M1 N$775 VI+ N$776 N$776 n_18_mm l=0.18u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M7 VO+ N$778 N$779 N$776 n_18_mm l=Ln w={{(Wncas/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wncas/1)}*5.4e-07)/2):(({(Wncas/1)}*4.9e-07+((1-1)*{(Wncas/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wncas/1)}*4.9e-07+(1-2)/2*({(Wncas/1)}*5.4e-07))/1):(({(Wncas/1)}*4.9e-07+((1-1)*{(Wncas/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wncas/1)}+5.4e-07):((2*({(Wncas/1)}+4.9e-07)+(1-1)*({(Wncas/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wncas/1)}+4.9e-07)+(1-2)*({(Wncas/1)}+5.4e-07))/1):((2*({(Wncas/1)}+4.9e-07)+(1-1)*({(Wncas/1)}+5.4e-07))/1))}
+  m=1
        E4 VO GROUND VO- VO+ 1
*
.end
