*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Thu Oct 24 2013 at 17:28:26

*
* Globals.
*
.global GROUND


*
* Component pathname : $MGC_DESIGN_KIT/symbols/MIMCAPS_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/MIMCAPS_MM/mimcaps_mm

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/OTA_SC1
*
        M16 VB2 VB2 VDD VDD p_18_mm l=Lin w={{({10*Win}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({10*Win}/1)}*5.4e-07)/2):(({({10*Win}/1)}*4.9e-07+((1-1)*{({10*Win}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({10*Win}/1)}*4.9e-07+(1-2)/2*({({10*Win}/1)}*5.4e-07))/1):(({({10*Win}/1)}*4.9e-07+((1-1)*{({10*Win}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({10*Win}/1)}+5.4e-07):((2*({({10*Win}/1)}+4.9e-07)+(1-1)*({({10*Win}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({10*Win}/1)}+4.9e-07)+(1-2)*({({10*Win}/1)}+5.4e-07))/1):((2*({({10*Win}/1)}+4.9e-07)+(1-1)*({({10*Win}/1)}+5.4e-07))/1))}
+  m=1
        I2 VB2 VB DC 100u
        M5 VOUT- N$598 VDD VDD p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M8 VOUT+ N$600 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M7 N$600 VCMFB GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        V3 N$338 GROUND PULSE ( 0V 1V 10nS 1nS 1nS 20nS 50nS )
        M4 VOUT+ N$548 VDD VDD p_18_mm l=Lp w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        C4 N$601 VOUT- Cc
        C3 VOUT+ N$600 Cc
        M2 N$600 VIN+ N$685 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        M6 N$601 VCMFB GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        X_S2D1 N$698 N$699 N$337 N$338 GROUND S2D
        V4 N$573 GROUND DC 0.9V
        E4 VCMFB GROUND N$572 N$573 -2
        M9 VOUT- N$601 GROUND GROUND n_18_mm l=Ln w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        C8 VIN- VOUT+ 200f
        C7 VIN+ VOUT- 200f
        C6 N$699 VIN- 200f
        C5 N$698 VIN+ 200f
        V2 N$337 GROUND DC 0.8V
        V1 VDD GROUND DC 1.8V
        E1 VO GROUND VOUT- VOUT+ -1
        M1 N$685 VB1 VDD VDD p_18_mm l=Lt w={{(Wt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wt/1)}*5.4e-07)/2):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wt/1)}*4.9e-07+(1-2)/2*({(Wt/1)}*5.4e-07))/1):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wt/1)}+5.4e-07):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wt/1)}+4.9e-07)+(1-2)*({(Wt/1)}+5.4e-07))/1):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  m=1
        E2 N$572 N$570 Vout+ 0 0.5
        M17 VB VB GROUND GROUND n_18_mm l=Ll w={{(Wl/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wl/1)}*5.4e-07)/2):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wl/1)}*4.9e-07+(1-2)/2*({(Wl/1)}*5.4e-07))/1):(({(Wl/1)}*4.9e-07+((1-1)*{(Wl/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wl/1)}+5.4e-07):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wl/1)}+4.9e-07)+(1-2)*({(Wl/1)}+5.4e-07))/1):((2*({(Wl/1)}+4.9e-07)+(1-1)*({(Wl/1)}+5.4e-07))/1))}
+  m=1
        I1 VB1 GROUND DC Ib
        E3 N$570 GROUND Vout- 0 0.5
        M12 VB1 VB1 VDD VDD p_18_mm l=Lt w={{(Wt/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wt/1)}*5.4e-07)/2):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wt/1)}*4.9e-07+(1-2)/2*({(Wt/1)}*5.4e-07))/1):(({(Wt/1)}*4.9e-07+((1-1)*{(Wt/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wt/1)}+5.4e-07):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wt/1)}+4.9e-07)+(1-2)*({(Wt/1)}+5.4e-07))/1):((2*({(Wt/1)}+4.9e-07)+(1-1)*({(Wt/1)}+5.4e-07))/1))}
+  m=1
        R1 N$548 VB1 40K
        XC2 N$598 N$601 mimcaps_mm w=Wc l=Lc m=1
        R2 VB1 N$598 40K
        M3 N$601 VIN- N$685 VDD p_18_mm l=Lin w={{(Win/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win/1)}*5.4e-07)/2):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win/1)}*4.9e-07+(1-2)/2*({(Win/1)}*5.4e-07))/1):(({(Win/1)}*4.9e-07+((1-1)*{(Win/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win/1)}+5.4e-07):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win/1)}+4.9e-07)+(1-2)*({(Win/1)}+5.4e-07))/1):((2*({(Win/1)}+4.9e-07)+(1-1)*({(Win/1)}+5.4e-07))/1))}
+  m=1
        XC1 N$548 N$600 mimcaps_mm w=Wc l=Lc m=1
*
.end
