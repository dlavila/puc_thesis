*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Tue Oct 29 2013 at 10:38:52

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/Tel_OTA_ideal
*
        V2 N$151 GROUND DC 0.9
        X_S2D1 VI+ VI- N$151 N$152 GROUND S2D
        M27 N$148 N$117 VDD2 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M26 N$117 N$113 N$148 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M25 N$117 N$99 N$147 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        C1 VO GROUND 2P
        I2 N$4 GROUND DC 300uA
        M23 VCASP N$113 VDD2 VDD2 p_18_mm l=2.2u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M22 N$113 N$113 VCASP VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M21 N$113 N$99 N$146 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M20 N$146 N$101 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M19 N$145 N$101 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M18 N$101 N$99 N$145 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M17 VCASN N$99 GROUND GROUND n_18_mm l=2.2u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M16 N$101 N$168 N$144 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M15 N$144 N$184 VDD2 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M10 N$168 N$168 N$184 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M13 N$78 N$184 VDD2 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M12 N$99 N$168 N$78 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M11 N$184 N$184 VDD2 VDD2 p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M14 N$99 N$99 VCASN GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        I1 N$168 VB4 DC 150uA
        V4 VDD2 GROUND DC 1.8V
        M24 N$147 N$101 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M28 VB4 VB4 GROUND GROUND n_18_mm l=0.45u w={{({Wn/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/2}/1)}*5.4e-07)/2):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/2}/1)}*4.9e-07+(1-2)/2*({({Wn/2}/1)}*5.4e-07))/1):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/2}/1)}+5.4e-07):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/2}/1)}+4.9e-07)+(1-2)*({({Wn/2}/1)}+5.4e-07))/1):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  m=1
        E1 N$56 GROUND VCASP N$55 250
        M9 N$54 N$7 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M8 N$55 N$7 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M7 N$7 N$57 N$54 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M6 VO N$56 N$55 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        E2 N$57 GROUND VCASP N$54 250
        E3 N$61 GROUND VCASN N$62 250
        E4 N$22 GROUND VCASN N$63 250
        M4 VO N$61 N$62 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M3 N$7 N$22 N$63 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M2 N$62 VI- N$4 GROUND n_18_mm l=0.18u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M1 N$63 VI+ N$4 GROUND n_18_mm l=0.18u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        V3 VDD GROUND DC 1.8V
        V1 N$152 GROUND DC 0V AC 1 0
*
.end
