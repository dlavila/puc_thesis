* Component: $LS_BUFFER/default.group/logic.views/NEW_BUFFER  Viewpoint: eldonet
.INCLUDE $LS_BUFFER/default.group/logic.views/NEW_BUFFER/eldonet/NEW_BUFFER_eldonet.spi
.INCLUDE $MGC_DESIGN_KIT/models/ELDO/include_all
.PROBE VX




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 
.PARAM Ln=0.45u 
.PARAM Lp=0.18u 
.PARAM Wn=40u 
.PARAM Wp=30u 
.PARAM Ib=10u 

.OPTION PROBOP2
.OPTION PROBOPX
.OP
.TRAN  0 100N 0 10p
