*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Mon Oct 28 2013 at 20:09:39

*
* Globals.
*
.global GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCP
*
.subckt AUX_FCP  VO VB1 VB2 VB3 VB4 VDD VI+ VI- VSS

        M6 N$252 VB1 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M15 VO VB2 N$248 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M14 N$249 VB2 N$246 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M13 N$246 N$249 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M19 N$248 N$249 VDD VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M30 N$251 VI- N$252 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M20 VO VB3 N$251 VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M21 N$251 VB4 VSS VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M17 N$249 VB3 N$253 VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
        M3 N$253 VI+ N$252 VDD p_18_mm l=0.45u w=1u ad=0.27p as=0.38p pd=1.54u
+  ps=2.26u m=4
        M10 N$253 VB4 VSS VSS n_18_mm l=0.45u w=0.5u ad=0.135p as=0.245p
+  pd=1.04u ps=1.98u m=2
.ends AUX_FCP

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCP_Bias
*
.subckt AUX_FCP_BIAS  VB1 VB2 VB3 VB4 IIN VDD VSS

        M12 VB1 VB3 N$32 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M7 N$32 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M4 N$31 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M2 VB2 VB3 N$31 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M1 VB2 VB2 N$33 VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M11 N$30 VB4 VSS VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M8 VB4 VB3 N$30 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M5 N$29 VB3 VSS VSS n_18_mm l=2.5u w=0.24u ad=0.118p as=0.118p pd=1.46u
+  ps=1.46u m=1
        M9 VB3 VB3 N$29 VSS n_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M18 VB4 IIN N$25 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M16 N$25 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M25 N$24 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M24 VB3 IIN N$24 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M23 N$34 VB1 VDD VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M29 N$22 N$22 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M28 IIN IIN N$22 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M26 VB1 VB2 N$34 VDD p_18_mm l=0.45u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
        M22 N$33 VB2 VDD VDD p_18_mm l=2.5u w=1u ad=0.49p as=0.49p pd=2.98u
+  ps=2.98u m=1
.ends AUX_FCP_BIAS

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCN_Bias
*
.subckt AUX_FCN_BIAS  VB1 VB2 VB3 VB4 IIN VDD VSS

        M7 N$15 VB1 VDD VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M6 VB1 VB2 N$15 VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M5 VB2 VB2 N$14 VDD p_18_mm l=0.45u w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
        M3 N$14 VB2 VDD VDD p_18_mm l=2.5u w=0.24u ad=0.118p as=0.118p pd=1.46u
+  ps=1.46u m=1
        M22 N$16 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M12 N$13 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M11 VB4 VB3 N$13 VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M9 N$12 VB3 VSS VSS n_18_mm l=2.5u w=0.75u ad=0.368p as=0.368p pd=2.48u
+  ps=2.48u m=1
        M8 VB3 VB3 N$12 VSS n_18_mm l=0.45u w=0.75u ad=0.368p as=0.368p
+  pd=2.48u ps=2.48u m=1
        M18 VB4 IIN N$11 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M16 N$11 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M25 N$10 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M24 VB3 IIN N$10 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p
+  pd=3.38u ps=3.38u m=1
        M27 N$17 VB4 VSS VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M29 N$8 N$8 VDD VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p pd=3.38u
+  ps=3.38u m=1
        M28 IIN IIN N$8 VDD p_18_mm l=0.45u w=1.2u ad=0.588p as=0.588p pd=3.38u
+  ps=3.38u m=1
        M26 VB1 VB3 N$17 VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
        M23 VB2 VB3 N$16 VSS n_18_mm l=0.45u w=0.75u ad=0.203p as=0.368p
+  pd=1.29u ps=2.48u m=2
.ends AUX_FCN_BIAS

*
* Component pathname : $AnalogIP/default.group/logic.views/AUX_FCN
*
.subckt AUX_FCN  VO VB1 VB2 VB3 VB4 VDD VI+ VI- VSS

        M19 N$681 VB1 VDD VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M10 VO VB3 N$614 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M20 N$616 N$678 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M21 N$678 VB3 N$616 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M2 N$677 VI+ N$619 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M15 VO VB2 N$681 VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M17 N$614 N$678 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M13 N$677 VB1 VDD VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
        M4 N$619 VB4 VSS VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M1 N$681 VI- N$619 VSS n_18_mm l=0.45u w=1.5u ad=0.405p as=0.735p
+  pd=2.04u ps=3.98u m=2
        M14 N$678 VB2 N$677 VDD p_18_mm l=0.45u w=0.4u ad=0.196p as=0.196p
+  pd=1.78u ps=1.78u m=1
.ends AUX_FCN

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/testMiniOpamps
*
        C2 GROUND VO2 60f
        C1 VO GROUND 60f
        I2 IREF2 GROUND DC 4uA
        V1 N$27 GROUND DC 0V AC 1 0
        V2 N$25 GROUND DC 1V
        X_AUX_FCP1 VO N$8 N$6 N$4 N$2 VDD N$40 N$51 GROUND AUX_FCP
        X_S2D1 N$40 N$51 N$25 N$27 GROUND S2D
        I1 IREF GROUND DC 6uA
        V3 VDD GROUND DC 1.8V
        X_AUX_FCP_BIAS1 N$8 N$6 N$4 N$2 IREF VDD GROUND AUX_FCP_BIAS
        X_AUX_FCN_BIAS1 N$34 N$35 N$36 N$37 IREF2 VDD GROUND AUX_FCN_BIAS
        X_AUX_FCN1 VO2 N$34 N$35 N$36 N$37 VDD N$40 N$51 GROUND AUX_FCN
*
.end
