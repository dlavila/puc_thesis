* Component: $SC_filter/default.group/logic.views/BIAS  Viewpoint: eldonet
.INCLUDE $SC_filter/default.group/logic.views/BIAS/eldonet/BIAS_eldonet.spi
.INCLUDE $MGC_DESIGN_KIT/models/ELDO/include_all
.PROBE VX
.PROBE I
.PROBE ISUB




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 

.OPTION PROBOP2
.OPTION PROBOPX
.OP
.TRAN  0 2m
