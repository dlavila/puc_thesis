*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Mon Sep 23 2013 at 16:00:29

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $SCF/default.group/logic.views/test
*
.subckt TEST  OUT IN VDD_ESC1 VSS

        M2 OUT IN VSS VSS n_18_mm l=$Lin w=0.24u ad=0.118p as=0.118p pd=1.46u
+  ps=1.46u m=1
        M1 OUT IN VDD_ESC1 VDD_ESC1 p_18_mm l=$Lin w=0.24u ad=0.118p as=0.118p
+  pd=1.46u ps=1.46u m=1
.ends TEST

*
* MAIN CELL: Component pathname : $SCF/default.group/logic.views/testTest
*
        X_TEST1 N$16 VIN VDD GROUND TEST
        V1 VDD GROUND DC 1.8V
        V2 VIN GROUND PULSE ( 0V 1.8V 0.01uS 0.01uS 0.5uS 1uS )
*
.end
