*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Fri Nov 29 2013 at 15:12:17

*
* Globals.
*
.global GROUND


*
* Component pathname : $MGC_DESIGN_KIT/symbols/MIMCAPS_MM [ELDOSPICE]
*
*       .include /usr/local/mentor/UMC180PDK/symbols/MIMCAPS_MM/mimcaps_mm

*
* Component pathname : $SC_filter/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* MAIN CELL: Component pathname : $RR_BUFFER/default.group/logic.views/BUFFER
*
        I1 N$880 GROUND DC Ib
        M43 N$880 N$880 VDD VDD p_18_mm l=0.45u w=6u ad=2.94p as=2.94p pd=12.98u
+  ps=12.98u m=1
        M39 VNCAS VB2 N$509 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        V6 VICM GROUND DC Vicm
        M33 VPCAS VPCAS N$421 VDD p_18_mm l=0.45u w={{({Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp}/1)}*5.4e-07)/2):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp}/1)}*4.9e-07+(1-2)/2*({({Wp}/1)}*5.4e-07))/1):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp}/1)}+5.4e-07):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp}/1)}+4.9e-07)+(1-2)*({({Wp}/1)}+5.4e-07))/1):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  m=1
        M31 N$808 VB4 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M13 N$841 VPCAS N$845 VDD p_18_mm l=0.45u w={{({Wp/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/2}/1)}*5.4e-07)/2):(({({Wp/2}/1)}*4.9e-07+((1-1)*{({Wp/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/2}/1)}*4.9e-07+(1-2)/2*({({Wp/2}/1)}*5.4e-07))/1):(({({Wp/2}/1)}*4.9e-07+((1-1)*{({Wp/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/2}/1)}+5.4e-07):((2*({({Wp/2}/1)}+4.9e-07)+(1-1)*({({Wp/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/2}/1)}+4.9e-07)+(1-2)*({({Wp/2}/1)}+5.4e-07))/1):((2*({({Wp/2}/1)}+4.9e-07)+(1-1)*({({Wp/2}/1)}+5.4e-07))/1))}
+  m=1
        M19 N$297 N$297 N$710 VDD p_18_mm l=Lin_p w={{({4*Win_p}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({4*Win_p}/1)}*5.4e-07)/2):(({({4*Win_p}/1)}*4.9e-07+((1-1)*{({4*Win_p}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({4*Win_p}/1)}*4.9e-07+(1-2)/2*({({4*Win_p}/1)}*5.4e-07))/1):(({({4*Win_p}/1)}*4.9e-07+((1-1)*{({4*Win_p}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({4*Win_p}/1)}+5.4e-07):((2*({({4*Win_p}/1)}+4.9e-07)+(1-1)*({({4*Win_p}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({4*Win_p}/1)}+4.9e-07)+(1-2)*({({4*Win_p}/1)}+5.4e-07))/1):((2*({({4*Win_p}/1)}+4.9e-07)+(1-1)*({({4*Win_p}/1)}+5.4e-07))/1))}
+  m=1
        MOUTP VO N$598 VDD VDD p_18_mm l=0.45u w={{({10*Wp}/10)}} ad={eval((10/2-trunc(10/2)==0)?(({({10*Wp}/10)}*5.4e-07)/2):(({({10*Wp}/10)}*4.9e-07+((10-1)*{({10*Wp}/10)}*5.4e-07)/2)/10))}
+  as={eval((10/2-trunc(10/2)==0)?((2*{({10*Wp}/10)}*4.9e-07+(10-2)/2*({({10*Wp}/10)}*5.4e-07))/10):(({({10*Wp}/10)}*4.9e-07+((10-1)*{({10*Wp}/10)}*5.4e-07)/2)/10))}
+  pd={eval((10/2-trunc(10/2)==0)?({({10*Wp}/10)}+5.4e-07):((2*({({10*Wp}/10)}+4.9e-07)+(10-1)*({({10*Wp}/10)}+5.4e-07))/10))}
+  ps={eval((10/2-trunc(10/2)==0)?((4*({({10*Wp}/10)}+4.9e-07)+(10-2)*({({10*Wp}/10)}+5.4e-07))/10):((2*({({10*Wp}/10)}+4.9e-07)+(10-1)*({({10*Wp}/10)}+5.4e-07))/10))}
+  m=10
        M3 N$722 VB1 VDD VDD p_18_mm l=0.45u w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M40 N$509 VB1 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M8 N$845 VNCAS N$841 GROUND n_18_mm l=0.45u w={{({Wn/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/2}/1)}*5.4e-07)/2):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/2}/1)}*4.9e-07+(1-2)/2*({({Wn/2}/1)}*5.4e-07))/1):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/2}/1)}+5.4e-07):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/2}/1)}+4.9e-07)+(1-2)*({({Wn/2}/1)}+5.4e-07))/1):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  m=1
        M42 VB3 N$880 VDD VDD p_18_mm l=0.45u w=6u ad=2.94p as=2.94p pd=12.98u
+  ps=12.98u m=1
        R1 N$598 N$868 Rr
        M37 N$810 VB1 VDD VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M27 N$805 VB4 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M23 VB4 VB3 N$511 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M12 N$598 VB2 N$854 VDD p_18_mm l=0.45u w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M38 VB1 VB2 N$810 VDD p_18_mm l=0.45u w={{(Wp/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wp/1)}*5.4e-07)/2):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wp/1)}*4.9e-07+(1-2)/2*({(Wp/1)}*5.4e-07))/1):(({(Wp/1)}*4.9e-07+((1-1)*{(Wp/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wp/1)}+5.4e-07):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wp/1)}+4.9e-07)+(1-2)*({(Wp/1)}+5.4e-07))/1):((2*({(Wp/1)}+4.9e-07)+(1-1)*({(Wp/1)}+5.4e-07))/1))}
+  m=1
        M21 VB3 VB3 N$793 GROUND n_18_mm l=0.45u w={{({Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn}/1)}*5.4e-07)/2):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn}/1)}*4.9e-07+(1-2)/2*({({Wn}/1)}*5.4e-07))/1):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn}/1)}+5.4e-07):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn}/1)}+4.9e-07)+(1-2)*({({Wn}/1)}+5.4e-07))/1):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  m=1
        M16 N$853 N$841 GROUND GROUND n_18_mm l=0.45u w={{({Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn}/1)}*5.4e-07)/2):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn}/1)}*4.9e-07+(1-2)/2*({({Wn}/1)}*5.4e-07))/1):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn}/1)}+5.4e-07):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn}/1)}+4.9e-07)+(1-2)*({({Wn}/1)}+5.4e-07))/1):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  m=1
        M20 N$297 N$297 N$709 GROUND n_18_mm l=Lin_n w={{({4*Win_n}/1)}}
+  ad={eval((1/2-trunc(1/2)==0)?(({({4*Win_n}/1)}*5.4e-07)/2):(({({4*Win_n}/1)}*4.9e-07+((1-1)*{({4*Win_n}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({4*Win_n}/1)}*4.9e-07+(1-2)/2*({({4*Win_n}/1)}*5.4e-07))/1):(({({4*Win_n}/1)}*4.9e-07+((1-1)*{({4*Win_n}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({4*Win_n}/1)}+5.4e-07):((2*({({4*Win_n}/1)}+4.9e-07)+(1-1)*({({4*Win_n}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({4*Win_n}/1)}+4.9e-07)+(1-2)*({({4*Win_n}/1)}+5.4e-07))/1):((2*({({4*Win_n}/1)}+4.9e-07)+(1-1)*({({4*Win_n}/1)}+5.4e-07))/1))}
+  m=1
        M35 N$482 N$482 GROUND GROUND n_18_mm l=0.45u w={{({2*Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wn}/1)}*5.4e-07)/2):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wn}/1)}*4.9e-07+(1-2)/2*({({2*Wn}/1)}*5.4e-07))/1):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wn}/1)}+5.4e-07):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wn}/1)}+4.9e-07)+(1-2)*({({2*Wn}/1)}+5.4e-07))/1):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  m=1
        M24 N$793 VB3 GROUND GROUND n_18_mm l=2.25u w={{({Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn}/1)}*5.4e-07)/2):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn}/1)}*4.9e-07+(1-2)/2*({({Wn}/1)}*5.4e-07))/1):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn}/1)}+5.4e-07):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn}/1)}+4.9e-07)+(1-2)*({({Wn}/1)}+5.4e-07))/1):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  m=1
        M10 N$845 VB2 N$844 VDD p_18_mm l=0.45u w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M34 N$421 N$421 VDD VDD p_18_mm l=0.45u w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M36 N$791 VB2 VDD VDD p_18_mm l=2.25u w={{({Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp}/1)}*5.4e-07)/2):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp}/1)}*4.9e-07+(1-2)/2*({({Wp}/1)}*5.4e-07))/1):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp}/1)}+5.4e-07):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp}/1)}+4.9e-07)+(1-2)*({({Wp}/1)}+5.4e-07))/1):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  m=1
        M4 N$709 VB3 N$725 GROUND n_18_mm l=0.45u w={{({2*Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wn}/1)}*5.4e-07)/2):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wn}/1)}*4.9e-07+(1-2)/2*({({2*Wn}/1)}*5.4e-07))/1):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wn}/1)}+5.4e-07):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wn}/1)}+4.9e-07)+(1-2)*({({2*Wn}/1)}+5.4e-07))/1):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  m=1
        M28 N$806 VB4 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M29 VB2 VB3 N$806 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        MIP2 N$853 VI+ N$710 VDD p_18_mm l=Lin_p w={{(Win_p/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win_p/1)}*5.4e-07)/2):(({(Win_p/1)}*4.9e-07+((1-1)*{(Win_p/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win_p/1)}*4.9e-07+(1-2)/2*({(Win_p/1)}*5.4e-07))/1):(({(Win_p/1)}*4.9e-07+((1-1)*{(Win_p/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win_p/1)}+5.4e-07):((2*({(Win_p/1)}+4.9e-07)+(1-1)*({(Win_p/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win_p/1)}+4.9e-07)+(1-2)*({(Win_p/1)}+5.4e-07))/1):((2*({(Win_p/1)}+4.9e-07)+(1-1)*({(Win_p/1)}+5.4e-07))/1))}
+  m=1
        M2 N$725 VB4 GROUND GROUND n_18_mm l=0.45u w={{({2*Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wn}/1)}*5.4e-07)/2):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wn}/1)}*4.9e-07+(1-2)/2*({({2*Wn}/1)}*5.4e-07))/1):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wn}/1)}+5.4e-07):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wn}/1)}+4.9e-07)+(1-2)*({({2*Wn}/1)}+5.4e-07))/1):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  m=1
        M17 N$854 VI+ N$709 GROUND n_18_mm l=Lin_n w={{(Win_n/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win_n/1)}*5.4e-07)/2):(({(Win_n/1)}*4.9e-07+((1-1)*{(Win_n/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win_n/1)}*4.9e-07+(1-2)/2*({(Win_n/1)}*5.4e-07))/1):(({(Win_n/1)}*4.9e-07+((1-1)*{(Win_n/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win_n/1)}+5.4e-07):((2*({(Win_n/1)}+4.9e-07)+(1-1)*({(Win_n/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win_n/1)}+4.9e-07)+(1-2)*({(Win_n/1)}+5.4e-07))/1):((2*({(Win_n/1)}+4.9e-07)+(1-1)*({(Win_n/1)}+5.4e-07))/1))}
+  m=1
        V1 N$865 GROUND DC 0V AC 1 0
        X_S2D1 VI+ VI- VICM N$865 GROUND S2D
        M41 VB4 N$880 VDD VDD p_18_mm l=0.45u w=6u ad=2.94p as=2.94p pd=12.98u
+  ps=12.98u m=1
        M18 N$840 VI- N$710 VDD p_18_mm l=Lin_p w={{(Win_p/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win_p/1)}*5.4e-07)/2):(({(Win_p/1)}*4.9e-07+((1-1)*{(Win_p/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win_p/1)}*4.9e-07+(1-2)/2*({(Win_p/1)}*5.4e-07))/1):(({(Win_p/1)}*4.9e-07+((1-1)*{(Win_p/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win_p/1)}+5.4e-07):((2*({(Win_p/1)}+4.9e-07)+(1-1)*({(Win_p/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win_p/1)}+4.9e-07)+(1-2)*({(Win_p/1)}+5.4e-07))/1):((2*({(Win_p/1)}+4.9e-07)+(1-1)*({(Win_p/1)}+5.4e-07))/1))}
+  m=1
        M14 N$751 VPCAS N$598 VDD p_18_mm l=0.45u w={{({Wp/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp/2}/1)}*5.4e-07)/2):(({({Wp/2}/1)}*4.9e-07+((1-1)*{({Wp/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp/2}/1)}*4.9e-07+(1-2)/2*({({Wp/2}/1)}*5.4e-07))/1):(({({Wp/2}/1)}*4.9e-07+((1-1)*{({Wp/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp/2}/1)}+5.4e-07):((2*({({Wp/2}/1)}+4.9e-07)+(1-1)*({({Wp/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp/2}/1)}+4.9e-07)+(1-2)*({({Wp/2}/1)}+5.4e-07))/1):((2*({({Wp/2}/1)}+4.9e-07)+(1-1)*({({Wp/2}/1)}+5.4e-07))/1))}
+  m=1
        V3 VDD GROUND DC 1.8V
        R2 N$751 N$870 Rr
        M32 VNCAS VNCAS N$482 GROUND n_18_mm l=0.45u w={{({Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn}/1)}*5.4e-07)/2):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn}/1)}*4.9e-07+(1-2)/2*({({Wn}/1)}*5.4e-07))/1):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn}/1)}+5.4e-07):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn}/1)}+4.9e-07)+(1-2)*({({Wn}/1)}+5.4e-07))/1):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  m=1
        M15 N$840 N$841 GROUND GROUND n_18_mm l=0.45u w={{({Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn}/1)}*5.4e-07)/2):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn}/1)}*4.9e-07+(1-2)/2*({({Wn}/1)}*5.4e-07))/1):(({({Wn}/1)}*4.9e-07+((1-1)*{({Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn}/1)}+5.4e-07):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn}/1)}+4.9e-07)+(1-2)*({({Wn}/1)}+5.4e-07))/1):((2*({({Wn}/1)}+4.9e-07)+(1-1)*({({Wn}/1)}+5.4e-07))/1))}
+  m=1
        M22 VB2 VB2 N$791 VDD p_18_mm l=0.45u w={{({Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp}/1)}*5.4e-07)/2):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp}/1)}*4.9e-07+(1-2)/2*({({Wp}/1)}*5.4e-07))/1):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp}/1)}+5.4e-07):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp}/1)}+4.9e-07)+(1-2)*({({Wp}/1)}+5.4e-07))/1):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  m=1
        M9 N$751 VB3 N$853 GROUND n_18_mm l=0.45u w={{({2*Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wn}/1)}*5.4e-07)/2):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wn}/1)}*4.9e-07+(1-2)/2*({({2*Wn}/1)}*5.4e-07))/1):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wn}/1)}+5.4e-07):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wn}/1)}+4.9e-07)+(1-2)*({({2*Wn}/1)}+5.4e-07))/1):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  m=1
        XC3 N$870 VO mimcaps_mm w=10u l=10u m=8
        XC2 N$868 VO mimcaps_mm w=10u l=10u m=8
        MOUTN VO N$751 GROUND GROUND n_18_mm l=0.45u w={{({10*Wn}/10)}}
+  ad={eval((10/2-trunc(10/2)==0)?(({({10*Wn}/10)}*5.4e-07)/2):(({({10*Wn}/10)}*4.9e-07+((10-1)*{({10*Wn}/10)}*5.4e-07)/2)/10))}
+  as={eval((10/2-trunc(10/2)==0)?((2*{({10*Wn}/10)}*4.9e-07+(10-2)/2*({({10*Wn}/10)}*5.4e-07))/10):(({({10*Wn}/10)}*4.9e-07+((10-1)*{({10*Wn}/10)}*5.4e-07)/2)/10))}
+  pd={eval((10/2-trunc(10/2)==0)?({({10*Wn}/10)}+5.4e-07):((2*({({10*Wn}/10)}+4.9e-07)+(10-1)*({({10*Wn}/10)}+5.4e-07))/10))}
+  ps={eval((10/2-trunc(10/2)==0)?((4*({({10*Wn}/10)}+4.9e-07)+(10-2)*({({10*Wn}/10)}+5.4e-07))/10):((2*({({10*Wn}/10)}+4.9e-07)+(10-1)*({({10*Wn}/10)}+5.4e-07))/10))}
+  m=10
        MIN1 N$844 VI- N$709 GROUND n_18_mm l=Lin_n w={{(Win_n/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Win_n/1)}*5.4e-07)/2):(({(Win_n/1)}*4.9e-07+((1-1)*{(Win_n/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Win_n/1)}*4.9e-07+(1-2)/2*({(Win_n/1)}*5.4e-07))/1):(({(Win_n/1)}*4.9e-07+((1-1)*{(Win_n/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Win_n/1)}+5.4e-07):((2*({(Win_n/1)}+4.9e-07)+(1-1)*({(Win_n/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Win_n/1)}+4.9e-07)+(1-2)*({(Win_n/1)}+5.4e-07))/1):((2*({(Win_n/1)}+4.9e-07)+(1-1)*({(Win_n/1)}+5.4e-07))/1))}
+  m=1
        M25 N$511 VB4 GROUND GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M30 VB1 VB3 N$808 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M1 N$710 VB2 N$722 VDD p_18_mm l=0.45u w={{({2*Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wp}/1)}*5.4e-07)/2):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wp}/1)}*4.9e-07+(1-2)/2*({({2*Wp}/1)}*5.4e-07))/1):(({({2*Wp}/1)}*4.9e-07+((1-1)*{({2*Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wp}/1)}+5.4e-07):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wp}/1)}+4.9e-07)+(1-2)*({({2*Wp}/1)}+5.4e-07))/1):((2*({({2*Wp}/1)}+4.9e-07)+(1-1)*({({2*Wp}/1)}+5.4e-07))/1))}
+  m=1
        M7 N$841 VB3 N$840 GROUND n_18_mm l=0.45u w={{({2*Wn}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({2*Wn}/1)}*5.4e-07)/2):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({2*Wn}/1)}*4.9e-07+(1-2)/2*({({2*Wn}/1)}*5.4e-07))/1):(({({2*Wn}/1)}*4.9e-07+((1-1)*{({2*Wn}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({2*Wn}/1)}+5.4e-07):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({2*Wn}/1)}+4.9e-07)+(1-2)*({({2*Wn}/1)}+5.4e-07))/1):((2*({({2*Wn}/1)}+4.9e-07)+(1-1)*({({2*Wn}/1)}+5.4e-07))/1))}
+  m=1
        C1 VO VICM 8P
        M26 VPCAS VB3 N$805 GROUND n_18_mm l=0.45u w={{(Wn/1)}} ad={eval((1/2-trunc(1/2)==0)?(({(Wn/1)}*5.4e-07)/2):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{(Wn/1)}*4.9e-07+(1-2)/2*({(Wn/1)}*5.4e-07))/1):(({(Wn/1)}*4.9e-07+((1-1)*{(Wn/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({(Wn/1)}+5.4e-07):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({(Wn/1)}+4.9e-07)+(1-2)*({(Wn/1)}+5.4e-07))/1):((2*({(Wn/1)}+4.9e-07)+(1-1)*({(Wn/1)}+5.4e-07))/1))}
+  m=1
        M6 N$854 N$845 VDD VDD p_18_mm l=0.45u w={{({Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp}/1)}*5.4e-07)/2):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp}/1)}*4.9e-07+(1-2)/2*({({Wp}/1)}*5.4e-07))/1):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp}/1)}+5.4e-07):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp}/1)}+4.9e-07)+(1-2)*({({Wp}/1)}+5.4e-07))/1):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  m=1
        M5 N$844 N$845 VDD VDD p_18_mm l=0.45u w={{({Wp}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wp}/1)}*5.4e-07)/2):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wp}/1)}*4.9e-07+(1-2)/2*({({Wp}/1)}*5.4e-07))/1):(({({Wp}/1)}*4.9e-07+((1-1)*{({Wp}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wp}/1)}+5.4e-07):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wp}/1)}+4.9e-07)+(1-2)*({({Wp}/1)}+5.4e-07))/1):((2*({({Wp}/1)}+4.9e-07)+(1-1)*({({Wp}/1)}+5.4e-07))/1))}
+  m=1
        M11 N$598 VNCAS N$751 GROUND n_18_mm l=0.45u w={{({Wn/2}/1)}} ad={eval((1/2-trunc(1/2)==0)?(({({Wn/2}/1)}*5.4e-07)/2):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  as={eval((1/2-trunc(1/2)==0)?((2*{({Wn/2}/1)}*4.9e-07+(1-2)/2*({({Wn/2}/1)}*5.4e-07))/1):(({({Wn/2}/1)}*4.9e-07+((1-1)*{({Wn/2}/1)}*5.4e-07)/2)/1))}
+  pd={eval((1/2-trunc(1/2)==0)?({({Wn/2}/1)}+5.4e-07):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  ps={eval((1/2-trunc(1/2)==0)?((4*({({Wn/2}/1)}+4.9e-07)+(1-2)*({({Wn/2}/1)}+5.4e-07))/1):((2*({({Wn/2}/1)}+4.9e-07)+(1-1)*({({Wn/2}/1)}+5.4e-07))/1))}
+  m=1
*
.end
