*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Tue Nov  5 2013 at 11:28:12

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $AnalogIP/default.group/logic.views/RFC_bias
*
.subckt RFC_BIAS  VB1 VB1T VB2 VB2T VB3 VB4 CURRENTIN VDD_ESC1 VSS

        M13 VB2T VB3 N$181 VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        M14 VB1T VB3 N$179 VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        M10 VB4 VB4 VSS VSS n_18_mm l=0.5u w=2u ad=0.98p as=0.98p pd=4.98u
+  ps=4.98u m=1
        M9 VB3 VB3 VB4 VSS n_18_mm l=0.18u w=2u ad=0.98p as=0.98p pd=4.98u
+  ps=4.98u m=1
        M4 VB3 CURRENTIN N$65 VDD_ESC1 p_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
        M18 N$181 VB4 VSS VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        M7 N$89 VB1T VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=0.5u ad=0.245p
+  as=0.245p pd=1.98u ps=1.98u m=1
        M21 VB2 VB3 N$175 VSS n_18_mm l=0.18u w=2u ad=0.98p as=0.98p pd=4.98u
+  ps=4.98u m=1
        M17 N$179 VB4 VSS VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        M12 VB1 VB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.5u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        M11 VB2 VB2 VB1 VDD_ESC1 p_18_mm l=0.18u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        MVB2 VB1T VB2T N$89 VDD_ESC1 p_18_mm l=0.18u w=0.5u ad=0.245p as=0.245p
+  pd=1.98u ps=1.98u m=1
        M1 VB2T VB2T N$91 VDD_ESC1 p_18_mm l=0.18u w=0.5u ad=0.245p as=0.245p
+  pd=1.98u ps=1.98u m=1
        M15 N$91 VB2T VDD_ESC1 VDD_ESC1 p_18_mm l=2u w=0.5u ad=0.245p as=0.245p
+  pd=1.98u ps=1.98u m=1
        M20 N$175 VB4 VSS VSS n_18_mm l=0.18u w=2u ad=0.98p as=0.98p pd=4.98u
+  ps=4.98u m=1
        M2 N$65 N$195 VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
        M5 CURRENTIN CURRENTIN N$195 VDD_ESC1 p_18_mm l=0.18u w=2u ad=0.98p
+  as=0.98p pd=4.98u ps=4.98u m=1
        M3 N$195 N$195 VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
.ends RFC_BIAS

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $AnalogIP/default.group/logic.views/RFC
*
.subckt RFC  VOUT+ VOUT- VB1 VB1T VB2 VB2T VB3 VB4 VDD_ESC1 VIN+ VIN- VOCM
+ VSS

        R2 N$727 N$336 1K
        R1 N$329 N$727 1K
        M13 N$669 VB4 VSS VSS n_18_mm l=0.5u w=16u ad=7.84p as=7.84p pd=32.98u
+  ps=32.98u m=1
        E3 N$336 VSS Vout- Vss 1
        M19 N$692 VB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.5u w=24u ad=11.76p as=11.76p
+  pd=48.98u ps=48.98u m=1
        E1 VDD_ESC1 CMFB1 N$727 VB1 -10
        M4 N$655 VB4 VSS VSS n_18_mm l=0.5u w=16u ad=7.84p as=7.84p pd=32.98u
+  ps=32.98u m=1
        M1A N$638 VIN+ N$718 VDD_ESC1 p_18_mm l=0.3u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M4B N$656 N$679 VSS VSS n_18_mm l=0.5u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M2 N$681 VB3 N$655 VSS n_18_mm l=0.18u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M0 N$717 VB1T VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=4u ad=1.96p as=1.96p
+  pd=8.98u ps=8.98u m=1
        M4A N$682 N$679 VSS VSS n_18_mm l=0.5u w=16u ad=7.84p as=7.84p pd=32.98u
+  ps=32.98u m=1
        M12 N$679 VB3 N$656 VSS n_18_mm l=0.18u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M5 VOUT- VB3 N$638 VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        M6 VOUT+ VB3 N$682 VSS n_18_mm l=0.18u w=8u ad=3.92p as=3.92p pd=16.98u
+  ps=16.98u m=1
        E2 N$329 VSS Vout+ Vss 1
        M9 N$692 CMFB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.5u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        M8 VOUT+ VB2 N$112 VDD_ESC1 p_18_mm l=0.18u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M10 N$112 CMFB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.5u w=8u ad=3.92p as=3.92p
+  pd=16.98u ps=16.98u m=1
        M18 N$682 VIN- N$718 VDD_ESC1 p_18_mm l=0.3u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M17 N$681 VIN- N$718 VDD_ESC1 p_18_mm l=0.3u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M16 N$679 VIN+ N$718 VDD_ESC1 p_18_mm l=0.3u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M11 N$681 VB3 N$653 VSS n_18_mm l=0.18u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M1 N$718 VB2T N$717 VDD_ESC1 p_18_mm l=0.18u w=4u ad=1.96p as=1.96p
+  pd=8.98u ps=8.98u m=1
        M3A N$638 N$681 VSS VSS n_18_mm l=0.5u w=16u ad=7.84p as=7.84p pd=32.98u
+  ps=32.98u m=1
        M3 N$679 VB3 N$669 VSS n_18_mm l=0.18u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M7 VOUT- VB2 N$692 VDD_ESC1 p_18_mm l=0.18u w=32u ad=15.68p as=15.68p
+  pd=64.98u ps=64.98u m=1
        M3B N$653 N$681 VSS VSS n_18_mm l=0.5u w=4u ad=1.96p as=1.96p pd=8.98u
+  ps=8.98u m=1
        M20 N$112 VB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.5u w=24u ad=11.76p as=11.76p
+  pd=48.98u ps=48.98u m=1
.ends RFC

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/testRFC
*
        C6 N$935 VO+ 1P
        C5 N$893 N$935 1P
        C4 N$931 VO- 1P
        C3 N$930 N$931 1P
        V2 N$331 GROUND DC Vicm
        I1 VDD N$659 DC 5u
        R4 GROUND VO- 10gig
        R3 VO+ GROUND 10gig
        V1 VDD GROUND DC 1.8V
        R2 VCM GROUND 1K
        E1 VO GROUND Vo+ Vo- 1
        R8 N$935 VO+ 10gig
        R7 N$893 N$935 10gig
        R6 N$931 VO- 10gig
        R5 N$930 N$931 10gig
        X_RFC_BIAS1 VB1 VB1T VB2 VB2T VB3 N$814 N$657 VDD GROUND RFC_BIAS
        M1 N$658 N$658 GROUND GROUND n_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
        V3 N$336 GROUND PULSE ( -0.1V 0.1V 10nS 1nS 1nS 20nS 50nS )
        C1 GROUND VO- 1P
        M4 N$657 N$659 N$660 GROUND n_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
        X_S2D1 N$930 N$893 N$331 N$336 GROUND S2D
        M2 N$660 N$658 GROUND GROUND n_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
        X_RFC1 VO- VO+ VB1 VB1T VB2 VB2T VB3 N$814 VDD N$935 N$931 VCM GROUND RFC
        C2 VO+ GROUND 1P
        R1 VDD VCM 1K
        M3 N$659 N$659 N$658 GROUND n_18_mm l=0.18u w=2u ad=0.98p as=0.98p
+  pd=4.98u ps=4.98u m=1
*
.end
