*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'dlavila' on Wed Oct  9 2013 at 14:00:02

*
* Globals.
*
.global GROUND VDD

*
* Component pathname : $AnalogIP/default.group/logic.views/s2d
*
.subckt S2D  VD+ VD- VICM VID VSS

        E3 N$2 VSS Vicm Vss 1
        E2 VD- N$2 Vss Vid 0.5
        E1 VD+ N$2 Vid Vss 0.5
.ends S2D

*
* Component pathname : $AnalogIP/default.group/logic.views/FFC
*
.subckt FFC  VO+ VO- VB1 VB2 VDD_ESC1 VI+ VI- VN VOCM VSS

        M11 N$179 VB2L N$83 VDD_ESC1 p_18_mm l=0.18u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        E1 CMFB VSS N$28 VOCM -20
        M19 VB2L VB2L VB1L VDD_ESC1 p_18_mm l=0.18u w=10u ad=2.7p as=3.14p
+  pd=10.54u ps=12.628u m=10
        M16 VB1L VB1L VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=6u ad=1.62p as=2.28p
+  pd=6.54u ps=9.76u m=4
        M0 N$202 VB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=10u ad=3.014p as=3.014p
+  pd=12.031u ps=12.031u m=7
        M13 VB2 VB2 VB1 VDD_ESC1 p_18_mm l=0.18u w=10u ad=3.014p as=3.014p
+  pd=12.031u ps=12.031u m=7
        M22 N$247 VB4 VSS VSS n_18_mm l=0.18u w=3u ad=1.47p as=1.47p pd=6.98u
+  ps=6.98u m=1
        M6 N$247 CMFB VSS VSS n_18_mm l=0.18u w=3u ad=1.03p as=1.03p pd=4.687u
+  ps=4.687u m=3
        M14 VO- N$188 N$238 VSS n_18_mm l=0.18u w=3u ad=0.81p as=1.14p pd=3.54u
+  ps=5.26u m=4
        M21 N$238 VB4 VSS VSS n_18_mm l=0.18u w=3u ad=1.47p as=1.47p pd=6.98u
+  ps=6.98u m=1
        M5 N$238 CMFB VSS VSS n_18_mm l=0.18u w=3u ad=1.03p as=1.03p pd=4.687u
+  ps=4.687u m=3
        M20 VB4 VB4 VSS VSS n_18_mm l=0.18u w=3u ad=0.81p as=1.14p pd=3.54u
+  ps=5.26u m=4
        M10 VSS VSS N$188 VDD_ESC1 p_18_mm l=0.18u w=0.6u ad=0.294p as=0.294p
+  pd=2.18u ps=2.18u m=1
        M12 VB1 VB1 VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=10u ad=3.014p as=3.014p
+  pd=12.031u ps=12.031u m=7
        I1 VB2 VB4 DC 700uA
        M1 N$238 VI+ N$34 VDD_ESC1 p_18_mm l=0.18u w=10u ad=2.7p as=3.14p
+  pd=10.54u ps=12.628u m=10
        M2 N$247 VI- N$34 VDD_ESC1 p_18_mm l=0.18u w=10u ad=2.7p as=3.14p
+  pd=10.54u ps=12.628u m=10
        M8 VO+ VB2L N$185 VDD_ESC1 p_18_mm l=0.18u w=10u ad=2.7p as=3.14p
+  pd=10.54u ps=12.628u m=10
        E2 N$28 N$30 Vout+ Vss 0.5
        E3 N$30 VSS Vout- Vss 0.5
        I2 VB2L VB4 DC 240uA
        M15 N$34 VB2 N$202 VDD_ESC1 p_18_mm l=0.18u w=10u ad=3.014p as=3.014p
+  pd=12.031u ps=12.031u m=7
        M3 N$83 VB1L VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=6u ad=1.62p as=2.28p
+  pd=6.54u ps=9.76u m=4
        M7 VO+ N$179 N$247 VSS n_18_mm l=0.18u w=3u ad=0.81p as=1.14p pd=3.54u
+  ps=5.26u m=4
        M17 N$185 VB1L VDD_ESC1 VDD_ESC1 p_18_mm l=0.18u w=6u ad=1.62p as=2.28p
+  pd=6.54u ps=9.76u m=4
        M4 VO- VB2L N$83 VDD_ESC1 p_18_mm l=0.18u w=10u ad=2.7p as=3.14p
+  pd=10.54u ps=12.628u m=10
        M9 N$188 VB2L N$185 VDD_ESC1 p_18_mm l=0.18u w=2.5u ad=1.225p as=1.225p
+  pd=5.98u ps=5.98u m=1
        M18 VSS VSS N$179 VDD_ESC1 p_18_mm l=0.18u w=0.6u ad=0.294p as=0.294p
+  pd=2.18u ps=2.18u m=1
.ends FFC

*
* MAIN CELL: Component pathname : $AnalogIP/default.group/logic.views/testFFC
*
        C2 N$30 GROUND 1P
        C1 GROUND N$31 1P
        V3 VDD GROUND DC 1.8V
        X_S2D1 N$22 N$15 N$8 N$9 GROUND S2D
        X_FFC1 N$30 N$31 N$21 N$20 VDD N$22 N$15 N$19 N$26 GROUND FFC
        V2 N$8 GROUND DC 1V
        V1 N$9 GROUND DC 0V AC 1 0
        E1 VO GROUND N$31 N$30 10
        V4 N$26 GROUND DC 0.9V
*
.end
